`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module picosoc_mem(
  input         clock,
  input         reset,
  input  [3:0]  wen,
  input  [21:0] addr,
  input  [31:0] wdata,
  output [31:0] rdata
);
  reg [31:0] mem_0;
  reg [31:0] _RAND_0;
  reg [31:0] mem_1;
  reg [31:0] _RAND_1;
  reg [31:0] mem_2;
  reg [31:0] _RAND_2;
  reg [31:0] mem_3;
  reg [31:0] _RAND_3;
  reg [31:0] mem_4;
  reg [31:0] _RAND_4;
  reg [31:0] mem_5;
  reg [31:0] _RAND_5;
  reg [31:0] mem_6;
  reg [31:0] _RAND_6;
  reg [31:0] mem_7;
  reg [31:0] _RAND_7;
  reg [31:0] mem_8;
  reg [31:0] _RAND_8;
  reg [31:0] mem_9;
  reg [31:0] _RAND_9;
  reg [31:0] mem_10;
  reg [31:0] _RAND_10;
  reg [31:0] mem_11;
  reg [31:0] _RAND_11;
  reg [31:0] mem_12;
  reg [31:0] _RAND_12;
  reg [31:0] mem_13;
  reg [31:0] _RAND_13;
  reg [31:0] mem_14;
  reg [31:0] _RAND_14;
  reg [31:0] mem_15;
  reg [31:0] _RAND_15;
  reg [31:0] mem_16;
  reg [31:0] _RAND_16;
  reg [31:0] mem_17;
  reg [31:0] _RAND_17;
  reg [31:0] mem_18;
  reg [31:0] _RAND_18;
  reg [31:0] mem_19;
  reg [31:0] _RAND_19;
  reg [31:0] mem_20;
  reg [31:0] _RAND_20;
  reg [31:0] mem_21;
  reg [31:0] _RAND_21;
  reg [31:0] mem_22;
  reg [31:0] _RAND_22;
  reg [31:0] mem_23;
  reg [31:0] _RAND_23;
  reg [31:0] mem_24;
  reg [31:0] _RAND_24;
  reg [31:0] mem_25;
  reg [31:0] _RAND_25;
  reg [31:0] mem_26;
  reg [31:0] _RAND_26;
  reg [31:0] mem_27;
  reg [31:0] _RAND_27;
  reg [31:0] mem_28;
  reg [31:0] _RAND_28;
  reg [31:0] mem_29;
  reg [31:0] _RAND_29;
  reg [31:0] mem_30;
  reg [31:0] _RAND_30;
  reg [31:0] mem_31;
  reg [31:0] _RAND_31;
  reg [31:0] mem_32;
  reg [31:0] _RAND_32;
  reg [31:0] mem_33;
  reg [31:0] _RAND_33;
  reg [31:0] mem_34;
  reg [31:0] _RAND_34;
  reg [31:0] mem_35;
  reg [31:0] _RAND_35;
  reg [31:0] mem_36;
  reg [31:0] _RAND_36;
  reg [31:0] mem_37;
  reg [31:0] _RAND_37;
  reg [31:0] mem_38;
  reg [31:0] _RAND_38;
  reg [31:0] mem_39;
  reg [31:0] _RAND_39;
  reg [31:0] mem_40;
  reg [31:0] _RAND_40;
  reg [31:0] mem_41;
  reg [31:0] _RAND_41;
  reg [31:0] mem_42;
  reg [31:0] _RAND_42;
  reg [31:0] mem_43;
  reg [31:0] _RAND_43;
  reg [31:0] mem_44;
  reg [31:0] _RAND_44;
  reg [31:0] mem_45;
  reg [31:0] _RAND_45;
  reg [31:0] mem_46;
  reg [31:0] _RAND_46;
  reg [31:0] mem_47;
  reg [31:0] _RAND_47;
  reg [31:0] mem_48;
  reg [31:0] _RAND_48;
  reg [31:0] mem_49;
  reg [31:0] _RAND_49;
  reg [31:0] mem_50;
  reg [31:0] _RAND_50;
  reg [31:0] mem_51;
  reg [31:0] _RAND_51;
  reg [31:0] mem_52;
  reg [31:0] _RAND_52;
  reg [31:0] mem_53;
  reg [31:0] _RAND_53;
  reg [31:0] mem_54;
  reg [31:0] _RAND_54;
  reg [31:0] mem_55;
  reg [31:0] _RAND_55;
  reg [31:0] mem_56;
  reg [31:0] _RAND_56;
  reg [31:0] mem_57;
  reg [31:0] _RAND_57;
  reg [31:0] mem_58;
  reg [31:0] _RAND_58;
  reg [31:0] mem_59;
  reg [31:0] _RAND_59;
  reg [31:0] mem_60;
  reg [31:0] _RAND_60;
  reg [31:0] mem_61;
  reg [31:0] _RAND_61;
  reg [31:0] mem_62;
  reg [31:0] _RAND_62;
  reg [31:0] mem_63;
  reg [31:0] _RAND_63;
  reg [31:0] mem_64;
  reg [31:0] _RAND_64;
  reg [31:0] mem_65;
  reg [31:0] _RAND_65;
  reg [31:0] mem_66;
  reg [31:0] _RAND_66;
  reg [31:0] mem_67;
  reg [31:0] _RAND_67;
  reg [31:0] mem_68;
  reg [31:0] _RAND_68;
  reg [31:0] mem_69;
  reg [31:0] _RAND_69;
  reg [31:0] mem_70;
  reg [31:0] _RAND_70;
  reg [31:0] mem_71;
  reg [31:0] _RAND_71;
  reg [31:0] mem_72;
  reg [31:0] _RAND_72;
  reg [31:0] mem_73;
  reg [31:0] _RAND_73;
  reg [31:0] mem_74;
  reg [31:0] _RAND_74;
  reg [31:0] mem_75;
  reg [31:0] _RAND_75;
  reg [31:0] mem_76;
  reg [31:0] _RAND_76;
  reg [31:0] mem_77;
  reg [31:0] _RAND_77;
  reg [31:0] mem_78;
  reg [31:0] _RAND_78;
  reg [31:0] mem_79;
  reg [31:0] _RAND_79;
  reg [31:0] mem_80;
  reg [31:0] _RAND_80;
  reg [31:0] mem_81;
  reg [31:0] _RAND_81;
  reg [31:0] mem_82;
  reg [31:0] _RAND_82;
  reg [31:0] mem_83;
  reg [31:0] _RAND_83;
  reg [31:0] mem_84;
  reg [31:0] _RAND_84;
  reg [31:0] mem_85;
  reg [31:0] _RAND_85;
  reg [31:0] mem_86;
  reg [31:0] _RAND_86;
  reg [31:0] mem_87;
  reg [31:0] _RAND_87;
  reg [31:0] mem_88;
  reg [31:0] _RAND_88;
  reg [31:0] mem_89;
  reg [31:0] _RAND_89;
  reg [31:0] mem_90;
  reg [31:0] _RAND_90;
  reg [31:0] mem_91;
  reg [31:0] _RAND_91;
  reg [31:0] mem_92;
  reg [31:0] _RAND_92;
  reg [31:0] mem_93;
  reg [31:0] _RAND_93;
  reg [31:0] mem_94;
  reg [31:0] _RAND_94;
  reg [31:0] mem_95;
  reg [31:0] _RAND_95;
  reg [31:0] mem_96;
  reg [31:0] _RAND_96;
  reg [31:0] mem_97;
  reg [31:0] _RAND_97;
  reg [31:0] mem_98;
  reg [31:0] _RAND_98;
  reg [31:0] mem_99;
  reg [31:0] _RAND_99;
  reg [31:0] mem_100;
  reg [31:0] _RAND_100;
  reg [31:0] mem_101;
  reg [31:0] _RAND_101;
  reg [31:0] mem_102;
  reg [31:0] _RAND_102;
  reg [31:0] mem_103;
  reg [31:0] _RAND_103;
  reg [31:0] mem_104;
  reg [31:0] _RAND_104;
  reg [31:0] mem_105;
  reg [31:0] _RAND_105;
  reg [31:0] mem_106;
  reg [31:0] _RAND_106;
  reg [31:0] mem_107;
  reg [31:0] _RAND_107;
  reg [31:0] mem_108;
  reg [31:0] _RAND_108;
  reg [31:0] mem_109;
  reg [31:0] _RAND_109;
  reg [31:0] mem_110;
  reg [31:0] _RAND_110;
  reg [31:0] mem_111;
  reg [31:0] _RAND_111;
  reg [31:0] mem_112;
  reg [31:0] _RAND_112;
  reg [31:0] mem_113;
  reg [31:0] _RAND_113;
  reg [31:0] mem_114;
  reg [31:0] _RAND_114;
  reg [31:0] mem_115;
  reg [31:0] _RAND_115;
  reg [31:0] mem_116;
  reg [31:0] _RAND_116;
  reg [31:0] mem_117;
  reg [31:0] _RAND_117;
  reg [31:0] mem_118;
  reg [31:0] _RAND_118;
  reg [31:0] mem_119;
  reg [31:0] _RAND_119;
  reg [31:0] mem_120;
  reg [31:0] _RAND_120;
  reg [31:0] mem_121;
  reg [31:0] _RAND_121;
  reg [31:0] mem_122;
  reg [31:0] _RAND_122;
  reg [31:0] mem_123;
  reg [31:0] _RAND_123;
  reg [31:0] mem_124;
  reg [31:0] _RAND_124;
  reg [31:0] mem_125;
  reg [31:0] _RAND_125;
  reg [31:0] mem_126;
  reg [31:0] _RAND_126;
  reg [31:0] mem_127;
  reg [31:0] _RAND_127;
  reg [31:0] mem_128;
  reg [31:0] _RAND_128;
  reg [31:0] mem_129;
  reg [31:0] _RAND_129;
  reg [31:0] mem_130;
  reg [31:0] _RAND_130;
  reg [31:0] mem_131;
  reg [31:0] _RAND_131;
  reg [31:0] mem_132;
  reg [31:0] _RAND_132;
  reg [31:0] mem_133;
  reg [31:0] _RAND_133;
  reg [31:0] mem_134;
  reg [31:0] _RAND_134;
  reg [31:0] mem_135;
  reg [31:0] _RAND_135;
  reg [31:0] mem_136;
  reg [31:0] _RAND_136;
  reg [31:0] mem_137;
  reg [31:0] _RAND_137;
  reg [31:0] mem_138;
  reg [31:0] _RAND_138;
  reg [31:0] mem_139;
  reg [31:0] _RAND_139;
  reg [31:0] mem_140;
  reg [31:0] _RAND_140;
  reg [31:0] mem_141;
  reg [31:0] _RAND_141;
  reg [31:0] mem_142;
  reg [31:0] _RAND_142;
  reg [31:0] mem_143;
  reg [31:0] _RAND_143;
  reg [31:0] mem_144;
  reg [31:0] _RAND_144;
  reg [31:0] mem_145;
  reg [31:0] _RAND_145;
  reg [31:0] mem_146;
  reg [31:0] _RAND_146;
  reg [31:0] mem_147;
  reg [31:0] _RAND_147;
  reg [31:0] mem_148;
  reg [31:0] _RAND_148;
  reg [31:0] mem_149;
  reg [31:0] _RAND_149;
  reg [31:0] mem_150;
  reg [31:0] _RAND_150;
  reg [31:0] mem_151;
  reg [31:0] _RAND_151;
  reg [31:0] mem_152;
  reg [31:0] _RAND_152;
  reg [31:0] mem_153;
  reg [31:0] _RAND_153;
  reg [31:0] mem_154;
  reg [31:0] _RAND_154;
  reg [31:0] mem_155;
  reg [31:0] _RAND_155;
  reg [31:0] mem_156;
  reg [31:0] _RAND_156;
  reg [31:0] mem_157;
  reg [31:0] _RAND_157;
  reg [31:0] mem_158;
  reg [31:0] _RAND_158;
  reg [31:0] mem_159;
  reg [31:0] _RAND_159;
  reg [31:0] mem_160;
  reg [31:0] _RAND_160;
  reg [31:0] mem_161;
  reg [31:0] _RAND_161;
  reg [31:0] mem_162;
  reg [31:0] _RAND_162;
  reg [31:0] mem_163;
  reg [31:0] _RAND_163;
  reg [31:0] mem_164;
  reg [31:0] _RAND_164;
  reg [31:0] mem_165;
  reg [31:0] _RAND_165;
  reg [31:0] mem_166;
  reg [31:0] _RAND_166;
  reg [31:0] mem_167;
  reg [31:0] _RAND_167;
  reg [31:0] mem_168;
  reg [31:0] _RAND_168;
  reg [31:0] mem_169;
  reg [31:0] _RAND_169;
  reg [31:0] mem_170;
  reg [31:0] _RAND_170;
  reg [31:0] mem_171;
  reg [31:0] _RAND_171;
  reg [31:0] mem_172;
  reg [31:0] _RAND_172;
  reg [31:0] mem_173;
  reg [31:0] _RAND_173;
  reg [31:0] mem_174;
  reg [31:0] _RAND_174;
  reg [31:0] mem_175;
  reg [31:0] _RAND_175;
  reg [31:0] mem_176;
  reg [31:0] _RAND_176;
  reg [31:0] mem_177;
  reg [31:0] _RAND_177;
  reg [31:0] mem_178;
  reg [31:0] _RAND_178;
  reg [31:0] mem_179;
  reg [31:0] _RAND_179;
  reg [31:0] mem_180;
  reg [31:0] _RAND_180;
  reg [31:0] mem_181;
  reg [31:0] _RAND_181;
  reg [31:0] mem_182;
  reg [31:0] _RAND_182;
  reg [31:0] mem_183;
  reg [31:0] _RAND_183;
  reg [31:0] mem_184;
  reg [31:0] _RAND_184;
  reg [31:0] mem_185;
  reg [31:0] _RAND_185;
  reg [31:0] mem_186;
  reg [31:0] _RAND_186;
  reg [31:0] mem_187;
  reg [31:0] _RAND_187;
  reg [31:0] mem_188;
  reg [31:0] _RAND_188;
  reg [31:0] mem_189;
  reg [31:0] _RAND_189;
  reg [31:0] mem_190;
  reg [31:0] _RAND_190;
  reg [31:0] mem_191;
  reg [31:0] _RAND_191;
  reg [31:0] mem_192;
  reg [31:0] _RAND_192;
  reg [31:0] mem_193;
  reg [31:0] _RAND_193;
  reg [31:0] mem_194;
  reg [31:0] _RAND_194;
  reg [31:0] mem_195;
  reg [31:0] _RAND_195;
  reg [31:0] mem_196;
  reg [31:0] _RAND_196;
  reg [31:0] mem_197;
  reg [31:0] _RAND_197;
  reg [31:0] mem_198;
  reg [31:0] _RAND_198;
  reg [31:0] mem_199;
  reg [31:0] _RAND_199;
  reg [31:0] mem_200;
  reg [31:0] _RAND_200;
  reg [31:0] mem_201;
  reg [31:0] _RAND_201;
  reg [31:0] mem_202;
  reg [31:0] _RAND_202;
  reg [31:0] mem_203;
  reg [31:0] _RAND_203;
  reg [31:0] mem_204;
  reg [31:0] _RAND_204;
  reg [31:0] mem_205;
  reg [31:0] _RAND_205;
  reg [31:0] mem_206;
  reg [31:0] _RAND_206;
  reg [31:0] mem_207;
  reg [31:0] _RAND_207;
  reg [31:0] mem_208;
  reg [31:0] _RAND_208;
  reg [31:0] mem_209;
  reg [31:0] _RAND_209;
  reg [31:0] mem_210;
  reg [31:0] _RAND_210;
  reg [31:0] mem_211;
  reg [31:0] _RAND_211;
  reg [31:0] mem_212;
  reg [31:0] _RAND_212;
  reg [31:0] mem_213;
  reg [31:0] _RAND_213;
  reg [31:0] mem_214;
  reg [31:0] _RAND_214;
  reg [31:0] mem_215;
  reg [31:0] _RAND_215;
  reg [31:0] mem_216;
  reg [31:0] _RAND_216;
  reg [31:0] mem_217;
  reg [31:0] _RAND_217;
  reg [31:0] mem_218;
  reg [31:0] _RAND_218;
  reg [31:0] mem_219;
  reg [31:0] _RAND_219;
  reg [31:0] mem_220;
  reg [31:0] _RAND_220;
  reg [31:0] mem_221;
  reg [31:0] _RAND_221;
  reg [31:0] mem_222;
  reg [31:0] _RAND_222;
  reg [31:0] mem_223;
  reg [31:0] _RAND_223;
  reg [31:0] mem_224;
  reg [31:0] _RAND_224;
  reg [31:0] mem_225;
  reg [31:0] _RAND_225;
  reg [31:0] mem_226;
  reg [31:0] _RAND_226;
  reg [31:0] mem_227;
  reg [31:0] _RAND_227;
  reg [31:0] mem_228;
  reg [31:0] _RAND_228;
  reg [31:0] mem_229;
  reg [31:0] _RAND_229;
  reg [31:0] mem_230;
  reg [31:0] _RAND_230;
  reg [31:0] mem_231;
  reg [31:0] _RAND_231;
  reg [31:0] mem_232;
  reg [31:0] _RAND_232;
  reg [31:0] mem_233;
  reg [31:0] _RAND_233;
  reg [31:0] mem_234;
  reg [31:0] _RAND_234;
  reg [31:0] mem_235;
  reg [31:0] _RAND_235;
  reg [31:0] mem_236;
  reg [31:0] _RAND_236;
  reg [31:0] mem_237;
  reg [31:0] _RAND_237;
  reg [31:0] mem_238;
  reg [31:0] _RAND_238;
  reg [31:0] mem_239;
  reg [31:0] _RAND_239;
  reg [31:0] mem_240;
  reg [31:0] _RAND_240;
  reg [31:0] mem_241;
  reg [31:0] _RAND_241;
  reg [31:0] mem_242;
  reg [31:0] _RAND_242;
  reg [31:0] mem_243;
  reg [31:0] _RAND_243;
  reg [31:0] mem_244;
  reg [31:0] _RAND_244;
  reg [31:0] mem_245;
  reg [31:0] _RAND_245;
  reg [31:0] mem_246;
  reg [31:0] _RAND_246;
  reg [31:0] mem_247;
  reg [31:0] _RAND_247;
  reg [31:0] mem_248;
  reg [31:0] _RAND_248;
  reg [31:0] mem_249;
  reg [31:0] _RAND_249;
  reg [31:0] mem_250;
  reg [31:0] _RAND_250;
  reg [31:0] mem_251;
  reg [31:0] _RAND_251;
  reg [31:0] mem_252;
  reg [31:0] _RAND_252;
  reg [31:0] mem_253;
  reg [31:0] _RAND_253;
  reg [31:0] mem_254;
  reg [31:0] _RAND_254;
  reg [31:0] mem_255;
  reg [31:0] _RAND_255;
  reg [31:0] mem_256;
  reg [31:0] _RAND_256;
  reg [31:0] mem_257;
  reg [31:0] _RAND_257;
  reg [31:0] mem_258;
  reg [31:0] _RAND_258;
  reg [31:0] mem_259;
  reg [31:0] _RAND_259;
  reg [31:0] mem_260;
  reg [31:0] _RAND_260;
  reg [31:0] mem_261;
  reg [31:0] _RAND_261;
  reg [31:0] mem_262;
  reg [31:0] _RAND_262;
  reg [31:0] mem_263;
  reg [31:0] _RAND_263;
  reg [31:0] mem_264;
  reg [31:0] _RAND_264;
  reg [31:0] mem_265;
  reg [31:0] _RAND_265;
  reg [31:0] mem_266;
  reg [31:0] _RAND_266;
  reg [31:0] mem_267;
  reg [31:0] _RAND_267;
  reg [31:0] mem_268;
  reg [31:0] _RAND_268;
  reg [31:0] mem_269;
  reg [31:0] _RAND_269;
  reg [31:0] mem_270;
  reg [31:0] _RAND_270;
  reg [31:0] mem_271;
  reg [31:0] _RAND_271;
  reg [31:0] mem_272;
  reg [31:0] _RAND_272;
  reg [31:0] mem_273;
  reg [31:0] _RAND_273;
  reg [31:0] mem_274;
  reg [31:0] _RAND_274;
  reg [31:0] mem_275;
  reg [31:0] _RAND_275;
  reg [31:0] mem_276;
  reg [31:0] _RAND_276;
  reg [31:0] mem_277;
  reg [31:0] _RAND_277;
  reg [31:0] mem_278;
  reg [31:0] _RAND_278;
  reg [31:0] mem_279;
  reg [31:0] _RAND_279;
  reg [31:0] mem_280;
  reg [31:0] _RAND_280;
  reg [31:0] mem_281;
  reg [31:0] _RAND_281;
  reg [31:0] mem_282;
  reg [31:0] _RAND_282;
  reg [31:0] mem_283;
  reg [31:0] _RAND_283;
  reg [31:0] mem_284;
  reg [31:0] _RAND_284;
  reg [31:0] mem_285;
  reg [31:0] _RAND_285;
  reg [31:0] mem_286;
  reg [31:0] _RAND_286;
  reg [31:0] mem_287;
  reg [31:0] _RAND_287;
  reg [31:0] mem_288;
  reg [31:0] _RAND_288;
  reg [31:0] mem_289;
  reg [31:0] _RAND_289;
  reg [31:0] mem_290;
  reg [31:0] _RAND_290;
  reg [31:0] mem_291;
  reg [31:0] _RAND_291;
  reg [31:0] mem_292;
  reg [31:0] _RAND_292;
  reg [31:0] mem_293;
  reg [31:0] _RAND_293;
  reg [31:0] mem_294;
  reg [31:0] _RAND_294;
  reg [31:0] mem_295;
  reg [31:0] _RAND_295;
  reg [31:0] mem_296;
  reg [31:0] _RAND_296;
  reg [31:0] mem_297;
  reg [31:0] _RAND_297;
  reg [31:0] mem_298;
  reg [31:0] _RAND_298;
  reg [31:0] mem_299;
  reg [31:0] _RAND_299;
  reg [31:0] mem_300;
  reg [31:0] _RAND_300;
  reg [31:0] mem_301;
  reg [31:0] _RAND_301;
  reg [31:0] mem_302;
  reg [31:0] _RAND_302;
  reg [31:0] mem_303;
  reg [31:0] _RAND_303;
  reg [31:0] mem_304;
  reg [31:0] _RAND_304;
  reg [31:0] mem_305;
  reg [31:0] _RAND_305;
  reg [31:0] mem_306;
  reg [31:0] _RAND_306;
  reg [31:0] mem_307;
  reg [31:0] _RAND_307;
  reg [31:0] mem_308;
  reg [31:0] _RAND_308;
  reg [31:0] mem_309;
  reg [31:0] _RAND_309;
  reg [31:0] mem_310;
  reg [31:0] _RAND_310;
  reg [31:0] mem_311;
  reg [31:0] _RAND_311;
  reg [31:0] mem_312;
  reg [31:0] _RAND_312;
  reg [31:0] mem_313;
  reg [31:0] _RAND_313;
  reg [31:0] mem_314;
  reg [31:0] _RAND_314;
  reg [31:0] mem_315;
  reg [31:0] _RAND_315;
  reg [31:0] mem_316;
  reg [31:0] _RAND_316;
  reg [31:0] mem_317;
  reg [31:0] _RAND_317;
  reg [31:0] mem_318;
  reg [31:0] _RAND_318;
  reg [31:0] mem_319;
  reg [31:0] _RAND_319;
  reg [31:0] mem_320;
  reg [31:0] _RAND_320;
  reg [31:0] mem_321;
  reg [31:0] _RAND_321;
  reg [31:0] mem_322;
  reg [31:0] _RAND_322;
  reg [31:0] mem_323;
  reg [31:0] _RAND_323;
  reg [31:0] mem_324;
  reg [31:0] _RAND_324;
  reg [31:0] mem_325;
  reg [31:0] _RAND_325;
  reg [31:0] mem_326;
  reg [31:0] _RAND_326;
  reg [31:0] mem_327;
  reg [31:0] _RAND_327;
  reg [31:0] mem_328;
  reg [31:0] _RAND_328;
  reg [31:0] mem_329;
  reg [31:0] _RAND_329;
  reg [31:0] mem_330;
  reg [31:0] _RAND_330;
  reg [31:0] mem_331;
  reg [31:0] _RAND_331;
  reg [31:0] mem_332;
  reg [31:0] _RAND_332;
  reg [31:0] mem_333;
  reg [31:0] _RAND_333;
  reg [31:0] mem_334;
  reg [31:0] _RAND_334;
  reg [31:0] mem_335;
  reg [31:0] _RAND_335;
  reg [31:0] mem_336;
  reg [31:0] _RAND_336;
  reg [31:0] mem_337;
  reg [31:0] _RAND_337;
  reg [31:0] mem_338;
  reg [31:0] _RAND_338;
  reg [31:0] mem_339;
  reg [31:0] _RAND_339;
  reg [31:0] mem_340;
  reg [31:0] _RAND_340;
  reg [31:0] mem_341;
  reg [31:0] _RAND_341;
  reg [31:0] mem_342;
  reg [31:0] _RAND_342;
  reg [31:0] mem_343;
  reg [31:0] _RAND_343;
  reg [31:0] mem_344;
  reg [31:0] _RAND_344;
  reg [31:0] mem_345;
  reg [31:0] _RAND_345;
  reg [31:0] mem_346;
  reg [31:0] _RAND_346;
  reg [31:0] mem_347;
  reg [31:0] _RAND_347;
  reg [31:0] mem_348;
  reg [31:0] _RAND_348;
  reg [31:0] mem_349;
  reg [31:0] _RAND_349;
  reg [31:0] mem_350;
  reg [31:0] _RAND_350;
  reg [31:0] mem_351;
  reg [31:0] _RAND_351;
  reg [31:0] mem_352;
  reg [31:0] _RAND_352;
  reg [31:0] mem_353;
  reg [31:0] _RAND_353;
  reg [31:0] mem_354;
  reg [31:0] _RAND_354;
  reg [31:0] mem_355;
  reg [31:0] _RAND_355;
  reg [31:0] mem_356;
  reg [31:0] _RAND_356;
  reg [31:0] mem_357;
  reg [31:0] _RAND_357;
  reg [31:0] mem_358;
  reg [31:0] _RAND_358;
  reg [31:0] mem_359;
  reg [31:0] _RAND_359;
  reg [31:0] mem_360;
  reg [31:0] _RAND_360;
  reg [31:0] mem_361;
  reg [31:0] _RAND_361;
  reg [31:0] mem_362;
  reg [31:0] _RAND_362;
  reg [31:0] mem_363;
  reg [31:0] _RAND_363;
  reg [31:0] mem_364;
  reg [31:0] _RAND_364;
  reg [31:0] mem_365;
  reg [31:0] _RAND_365;
  reg [31:0] mem_366;
  reg [31:0] _RAND_366;
  reg [31:0] mem_367;
  reg [31:0] _RAND_367;
  reg [31:0] mem_368;
  reg [31:0] _RAND_368;
  reg [31:0] mem_369;
  reg [31:0] _RAND_369;
  reg [31:0] mem_370;
  reg [31:0] _RAND_370;
  reg [31:0] mem_371;
  reg [31:0] _RAND_371;
  reg [31:0] mem_372;
  reg [31:0] _RAND_372;
  reg [31:0] mem_373;
  reg [31:0] _RAND_373;
  reg [31:0] mem_374;
  reg [31:0] _RAND_374;
  reg [31:0] mem_375;
  reg [31:0] _RAND_375;
  reg [31:0] mem_376;
  reg [31:0] _RAND_376;
  reg [31:0] mem_377;
  reg [31:0] _RAND_377;
  reg [31:0] mem_378;
  reg [31:0] _RAND_378;
  reg [31:0] mem_379;
  reg [31:0] _RAND_379;
  reg [31:0] mem_380;
  reg [31:0] _RAND_380;
  reg [31:0] mem_381;
  reg [31:0] _RAND_381;
  reg [31:0] mem_382;
  reg [31:0] _RAND_382;
  reg [31:0] mem_383;
  reg [31:0] _RAND_383;
  reg [31:0] mem_384;
  reg [31:0] _RAND_384;
  reg [31:0] mem_385;
  reg [31:0] _RAND_385;
  reg [31:0] mem_386;
  reg [31:0] _RAND_386;
  reg [31:0] mem_387;
  reg [31:0] _RAND_387;
  reg [31:0] mem_388;
  reg [31:0] _RAND_388;
  reg [31:0] mem_389;
  reg [31:0] _RAND_389;
  reg [31:0] mem_390;
  reg [31:0] _RAND_390;
  reg [31:0] mem_391;
  reg [31:0] _RAND_391;
  reg [31:0] mem_392;
  reg [31:0] _RAND_392;
  reg [31:0] mem_393;
  reg [31:0] _RAND_393;
  reg [31:0] mem_394;
  reg [31:0] _RAND_394;
  reg [31:0] mem_395;
  reg [31:0] _RAND_395;
  reg [31:0] mem_396;
  reg [31:0] _RAND_396;
  reg [31:0] mem_397;
  reg [31:0] _RAND_397;
  reg [31:0] mem_398;
  reg [31:0] _RAND_398;
  reg [31:0] mem_399;
  reg [31:0] _RAND_399;
  reg [31:0] mem_400;
  reg [31:0] _RAND_400;
  reg [31:0] mem_401;
  reg [31:0] _RAND_401;
  reg [31:0] mem_402;
  reg [31:0] _RAND_402;
  reg [31:0] mem_403;
  reg [31:0] _RAND_403;
  reg [31:0] mem_404;
  reg [31:0] _RAND_404;
  reg [31:0] mem_405;
  reg [31:0] _RAND_405;
  reg [31:0] mem_406;
  reg [31:0] _RAND_406;
  reg [31:0] mem_407;
  reg [31:0] _RAND_407;
  reg [31:0] mem_408;
  reg [31:0] _RAND_408;
  reg [31:0] mem_409;
  reg [31:0] _RAND_409;
  reg [31:0] mem_410;
  reg [31:0] _RAND_410;
  reg [31:0] mem_411;
  reg [31:0] _RAND_411;
  reg [31:0] mem_412;
  reg [31:0] _RAND_412;
  reg [31:0] mem_413;
  reg [31:0] _RAND_413;
  reg [31:0] mem_414;
  reg [31:0] _RAND_414;
  reg [31:0] mem_415;
  reg [31:0] _RAND_415;
  reg [31:0] mem_416;
  reg [31:0] _RAND_416;
  reg [31:0] mem_417;
  reg [31:0] _RAND_417;
  reg [31:0] mem_418;
  reg [31:0] _RAND_418;
  reg [31:0] mem_419;
  reg [31:0] _RAND_419;
  reg [31:0] mem_420;
  reg [31:0] _RAND_420;
  reg [31:0] mem_421;
  reg [31:0] _RAND_421;
  reg [31:0] mem_422;
  reg [31:0] _RAND_422;
  reg [31:0] mem_423;
  reg [31:0] _RAND_423;
  reg [31:0] mem_424;
  reg [31:0] _RAND_424;
  reg [31:0] mem_425;
  reg [31:0] _RAND_425;
  reg [31:0] mem_426;
  reg [31:0] _RAND_426;
  reg [31:0] mem_427;
  reg [31:0] _RAND_427;
  reg [31:0] mem_428;
  reg [31:0] _RAND_428;
  reg [31:0] mem_429;
  reg [31:0] _RAND_429;
  reg [31:0] mem_430;
  reg [31:0] _RAND_430;
  reg [31:0] mem_431;
  reg [31:0] _RAND_431;
  reg [31:0] mem_432;
  reg [31:0] _RAND_432;
  reg [31:0] mem_433;
  reg [31:0] _RAND_433;
  reg [31:0] mem_434;
  reg [31:0] _RAND_434;
  reg [31:0] mem_435;
  reg [31:0] _RAND_435;
  reg [31:0] mem_436;
  reg [31:0] _RAND_436;
  reg [31:0] mem_437;
  reg [31:0] _RAND_437;
  reg [31:0] mem_438;
  reg [31:0] _RAND_438;
  reg [31:0] mem_439;
  reg [31:0] _RAND_439;
  reg [31:0] mem_440;
  reg [31:0] _RAND_440;
  reg [31:0] mem_441;
  reg [31:0] _RAND_441;
  reg [31:0] mem_442;
  reg [31:0] _RAND_442;
  reg [31:0] mem_443;
  reg [31:0] _RAND_443;
  reg [31:0] mem_444;
  reg [31:0] _RAND_444;
  reg [31:0] mem_445;
  reg [31:0] _RAND_445;
  reg [31:0] mem_446;
  reg [31:0] _RAND_446;
  reg [31:0] mem_447;
  reg [31:0] _RAND_447;
  reg [31:0] mem_448;
  reg [31:0] _RAND_448;
  reg [31:0] mem_449;
  reg [31:0] _RAND_449;
  reg [31:0] mem_450;
  reg [31:0] _RAND_450;
  reg [31:0] mem_451;
  reg [31:0] _RAND_451;
  reg [31:0] mem_452;
  reg [31:0] _RAND_452;
  reg [31:0] mem_453;
  reg [31:0] _RAND_453;
  reg [31:0] mem_454;
  reg [31:0] _RAND_454;
  reg [31:0] mem_455;
  reg [31:0] _RAND_455;
  reg [31:0] mem_456;
  reg [31:0] _RAND_456;
  reg [31:0] mem_457;
  reg [31:0] _RAND_457;
  reg [31:0] mem_458;
  reg [31:0] _RAND_458;
  reg [31:0] mem_459;
  reg [31:0] _RAND_459;
  reg [31:0] mem_460;
  reg [31:0] _RAND_460;
  reg [31:0] mem_461;
  reg [31:0] _RAND_461;
  reg [31:0] mem_462;
  reg [31:0] _RAND_462;
  reg [31:0] mem_463;
  reg [31:0] _RAND_463;
  reg [31:0] mem_464;
  reg [31:0] _RAND_464;
  reg [31:0] mem_465;
  reg [31:0] _RAND_465;
  reg [31:0] mem_466;
  reg [31:0] _RAND_466;
  reg [31:0] mem_467;
  reg [31:0] _RAND_467;
  reg [31:0] mem_468;
  reg [31:0] _RAND_468;
  reg [31:0] mem_469;
  reg [31:0] _RAND_469;
  reg [31:0] mem_470;
  reg [31:0] _RAND_470;
  reg [31:0] mem_471;
  reg [31:0] _RAND_471;
  reg [31:0] mem_472;
  reg [31:0] _RAND_472;
  reg [31:0] mem_473;
  reg [31:0] _RAND_473;
  reg [31:0] mem_474;
  reg [31:0] _RAND_474;
  reg [31:0] mem_475;
  reg [31:0] _RAND_475;
  reg [31:0] mem_476;
  reg [31:0] _RAND_476;
  reg [31:0] mem_477;
  reg [31:0] _RAND_477;
  reg [31:0] mem_478;
  reg [31:0] _RAND_478;
  reg [31:0] mem_479;
  reg [31:0] _RAND_479;
  reg [31:0] mem_480;
  reg [31:0] _RAND_480;
  reg [31:0] mem_481;
  reg [31:0] _RAND_481;
  reg [31:0] mem_482;
  reg [31:0] _RAND_482;
  reg [31:0] mem_483;
  reg [31:0] _RAND_483;
  reg [31:0] mem_484;
  reg [31:0] _RAND_484;
  reg [31:0] mem_485;
  reg [31:0] _RAND_485;
  reg [31:0] mem_486;
  reg [31:0] _RAND_486;
  reg [31:0] mem_487;
  reg [31:0] _RAND_487;
  reg [31:0] mem_488;
  reg [31:0] _RAND_488;
  reg [31:0] mem_489;
  reg [31:0] _RAND_489;
  reg [31:0] mem_490;
  reg [31:0] _RAND_490;
  reg [31:0] mem_491;
  reg [31:0] _RAND_491;
  reg [31:0] mem_492;
  reg [31:0] _RAND_492;
  reg [31:0] mem_493;
  reg [31:0] _RAND_493;
  reg [31:0] mem_494;
  reg [31:0] _RAND_494;
  reg [31:0] mem_495;
  reg [31:0] _RAND_495;
  reg [31:0] mem_496;
  reg [31:0] _RAND_496;
  reg [31:0] mem_497;
  reg [31:0] _RAND_497;
  reg [31:0] mem_498;
  reg [31:0] _RAND_498;
  reg [31:0] mem_499;
  reg [31:0] _RAND_499;
  reg [31:0] mem_500;
  reg [31:0] _RAND_500;
  reg [31:0] mem_501;
  reg [31:0] _RAND_501;
  reg [31:0] mem_502;
  reg [31:0] _RAND_502;
  reg [31:0] mem_503;
  reg [31:0] _RAND_503;
  reg [31:0] mem_504;
  reg [31:0] _RAND_504;
  reg [31:0] mem_505;
  reg [31:0] _RAND_505;
  reg [31:0] mem_506;
  reg [31:0] _RAND_506;
  reg [31:0] mem_507;
  reg [31:0] _RAND_507;
  reg [31:0] mem_508;
  reg [31:0] _RAND_508;
  reg [31:0] mem_509;
  reg [31:0] _RAND_509;
  reg [31:0] mem_510;
  reg [31:0] _RAND_510;
  reg [31:0] mem_511;
  reg [31:0] _RAND_511;
  reg [31:0] mem_512;
  reg [31:0] _RAND_512;
  reg [31:0] mem_513;
  reg [31:0] _RAND_513;
  reg [31:0] mem_514;
  reg [31:0] _RAND_514;
  reg [31:0] mem_515;
  reg [31:0] _RAND_515;
  reg [31:0] mem_516;
  reg [31:0] _RAND_516;
  reg [31:0] mem_517;
  reg [31:0] _RAND_517;
  reg [31:0] mem_518;
  reg [31:0] _RAND_518;
  reg [31:0] mem_519;
  reg [31:0] _RAND_519;
  reg [31:0] mem_520;
  reg [31:0] _RAND_520;
  reg [31:0] mem_521;
  reg [31:0] _RAND_521;
  reg [31:0] mem_522;
  reg [31:0] _RAND_522;
  reg [31:0] mem_523;
  reg [31:0] _RAND_523;
  reg [31:0] mem_524;
  reg [31:0] _RAND_524;
  reg [31:0] mem_525;
  reg [31:0] _RAND_525;
  reg [31:0] mem_526;
  reg [31:0] _RAND_526;
  reg [31:0] mem_527;
  reg [31:0] _RAND_527;
  reg [31:0] mem_528;
  reg [31:0] _RAND_528;
  reg [31:0] mem_529;
  reg [31:0] _RAND_529;
  reg [31:0] mem_530;
  reg [31:0] _RAND_530;
  reg [31:0] mem_531;
  reg [31:0] _RAND_531;
  reg [31:0] mem_532;
  reg [31:0] _RAND_532;
  reg [31:0] mem_533;
  reg [31:0] _RAND_533;
  reg [31:0] mem_534;
  reg [31:0] _RAND_534;
  reg [31:0] mem_535;
  reg [31:0] _RAND_535;
  reg [31:0] mem_536;
  reg [31:0] _RAND_536;
  reg [31:0] mem_537;
  reg [31:0] _RAND_537;
  reg [31:0] mem_538;
  reg [31:0] _RAND_538;
  reg [31:0] mem_539;
  reg [31:0] _RAND_539;
  reg [31:0] mem_540;
  reg [31:0] _RAND_540;
  reg [31:0] mem_541;
  reg [31:0] _RAND_541;
  reg [31:0] mem_542;
  reg [31:0] _RAND_542;
  reg [31:0] mem_543;
  reg [31:0] _RAND_543;
  reg [31:0] mem_544;
  reg [31:0] _RAND_544;
  reg [31:0] mem_545;
  reg [31:0] _RAND_545;
  reg [31:0] mem_546;
  reg [31:0] _RAND_546;
  reg [31:0] mem_547;
  reg [31:0] _RAND_547;
  reg [31:0] mem_548;
  reg [31:0] _RAND_548;
  reg [31:0] mem_549;
  reg [31:0] _RAND_549;
  reg [31:0] mem_550;
  reg [31:0] _RAND_550;
  reg [31:0] mem_551;
  reg [31:0] _RAND_551;
  reg [31:0] mem_552;
  reg [31:0] _RAND_552;
  reg [31:0] mem_553;
  reg [31:0] _RAND_553;
  reg [31:0] mem_554;
  reg [31:0] _RAND_554;
  reg [31:0] mem_555;
  reg [31:0] _RAND_555;
  reg [31:0] mem_556;
  reg [31:0] _RAND_556;
  reg [31:0] mem_557;
  reg [31:0] _RAND_557;
  reg [31:0] mem_558;
  reg [31:0] _RAND_558;
  reg [31:0] mem_559;
  reg [31:0] _RAND_559;
  reg [31:0] mem_560;
  reg [31:0] _RAND_560;
  reg [31:0] mem_561;
  reg [31:0] _RAND_561;
  reg [31:0] mem_562;
  reg [31:0] _RAND_562;
  reg [31:0] mem_563;
  reg [31:0] _RAND_563;
  reg [31:0] mem_564;
  reg [31:0] _RAND_564;
  reg [31:0] mem_565;
  reg [31:0] _RAND_565;
  reg [31:0] mem_566;
  reg [31:0] _RAND_566;
  reg [31:0] mem_567;
  reg [31:0] _RAND_567;
  reg [31:0] mem_568;
  reg [31:0] _RAND_568;
  reg [31:0] mem_569;
  reg [31:0] _RAND_569;
  reg [31:0] mem_570;
  reg [31:0] _RAND_570;
  reg [31:0] mem_571;
  reg [31:0] _RAND_571;
  reg [31:0] mem_572;
  reg [31:0] _RAND_572;
  reg [31:0] mem_573;
  reg [31:0] _RAND_573;
  reg [31:0] mem_574;
  reg [31:0] _RAND_574;
  reg [31:0] mem_575;
  reg [31:0] _RAND_575;
  reg [31:0] mem_576;
  reg [31:0] _RAND_576;
  reg [31:0] mem_577;
  reg [31:0] _RAND_577;
  reg [31:0] mem_578;
  reg [31:0] _RAND_578;
  reg [31:0] mem_579;
  reg [31:0] _RAND_579;
  reg [31:0] mem_580;
  reg [31:0] _RAND_580;
  reg [31:0] mem_581;
  reg [31:0] _RAND_581;
  reg [31:0] mem_582;
  reg [31:0] _RAND_582;
  reg [31:0] mem_583;
  reg [31:0] _RAND_583;
  reg [31:0] mem_584;
  reg [31:0] _RAND_584;
  reg [31:0] mem_585;
  reg [31:0] _RAND_585;
  reg [31:0] mem_586;
  reg [31:0] _RAND_586;
  reg [31:0] mem_587;
  reg [31:0] _RAND_587;
  reg [31:0] mem_588;
  reg [31:0] _RAND_588;
  reg [31:0] mem_589;
  reg [31:0] _RAND_589;
  reg [31:0] mem_590;
  reg [31:0] _RAND_590;
  reg [31:0] mem_591;
  reg [31:0] _RAND_591;
  reg [31:0] mem_592;
  reg [31:0] _RAND_592;
  reg [31:0] mem_593;
  reg [31:0] _RAND_593;
  reg [31:0] mem_594;
  reg [31:0] _RAND_594;
  reg [31:0] mem_595;
  reg [31:0] _RAND_595;
  reg [31:0] mem_596;
  reg [31:0] _RAND_596;
  reg [31:0] mem_597;
  reg [31:0] _RAND_597;
  reg [31:0] mem_598;
  reg [31:0] _RAND_598;
  reg [31:0] mem_599;
  reg [31:0] _RAND_599;
  reg [31:0] mem_600;
  reg [31:0] _RAND_600;
  reg [31:0] mem_601;
  reg [31:0] _RAND_601;
  reg [31:0] mem_602;
  reg [31:0] _RAND_602;
  reg [31:0] mem_603;
  reg [31:0] _RAND_603;
  reg [31:0] mem_604;
  reg [31:0] _RAND_604;
  reg [31:0] mem_605;
  reg [31:0] _RAND_605;
  reg [31:0] mem_606;
  reg [31:0] _RAND_606;
  reg [31:0] mem_607;
  reg [31:0] _RAND_607;
  reg [31:0] mem_608;
  reg [31:0] _RAND_608;
  reg [31:0] mem_609;
  reg [31:0] _RAND_609;
  reg [31:0] mem_610;
  reg [31:0] _RAND_610;
  reg [31:0] mem_611;
  reg [31:0] _RAND_611;
  reg [31:0] mem_612;
  reg [31:0] _RAND_612;
  reg [31:0] mem_613;
  reg [31:0] _RAND_613;
  reg [31:0] mem_614;
  reg [31:0] _RAND_614;
  reg [31:0] mem_615;
  reg [31:0] _RAND_615;
  reg [31:0] mem_616;
  reg [31:0] _RAND_616;
  reg [31:0] mem_617;
  reg [31:0] _RAND_617;
  reg [31:0] mem_618;
  reg [31:0] _RAND_618;
  reg [31:0] mem_619;
  reg [31:0] _RAND_619;
  reg [31:0] mem_620;
  reg [31:0] _RAND_620;
  reg [31:0] mem_621;
  reg [31:0] _RAND_621;
  reg [31:0] mem_622;
  reg [31:0] _RAND_622;
  reg [31:0] mem_623;
  reg [31:0] _RAND_623;
  reg [31:0] mem_624;
  reg [31:0] _RAND_624;
  reg [31:0] mem_625;
  reg [31:0] _RAND_625;
  reg [31:0] mem_626;
  reg [31:0] _RAND_626;
  reg [31:0] mem_627;
  reg [31:0] _RAND_627;
  reg [31:0] mem_628;
  reg [31:0] _RAND_628;
  reg [31:0] mem_629;
  reg [31:0] _RAND_629;
  reg [31:0] mem_630;
  reg [31:0] _RAND_630;
  reg [31:0] mem_631;
  reg [31:0] _RAND_631;
  reg [31:0] mem_632;
  reg [31:0] _RAND_632;
  reg [31:0] mem_633;
  reg [31:0] _RAND_633;
  reg [31:0] mem_634;
  reg [31:0] _RAND_634;
  reg [31:0] mem_635;
  reg [31:0] _RAND_635;
  reg [31:0] mem_636;
  reg [31:0] _RAND_636;
  reg [31:0] mem_637;
  reg [31:0] _RAND_637;
  reg [31:0] mem_638;
  reg [31:0] _RAND_638;
  reg [31:0] mem_639;
  reg [31:0] _RAND_639;
  reg [31:0] mem_640;
  reg [31:0] _RAND_640;
  reg [31:0] mem_641;
  reg [31:0] _RAND_641;
  reg [31:0] mem_642;
  reg [31:0] _RAND_642;
  reg [31:0] mem_643;
  reg [31:0] _RAND_643;
  reg [31:0] mem_644;
  reg [31:0] _RAND_644;
  reg [31:0] mem_645;
  reg [31:0] _RAND_645;
  reg [31:0] mem_646;
  reg [31:0] _RAND_646;
  reg [31:0] mem_647;
  reg [31:0] _RAND_647;
  reg [31:0] mem_648;
  reg [31:0] _RAND_648;
  reg [31:0] mem_649;
  reg [31:0] _RAND_649;
  reg [31:0] mem_650;
  reg [31:0] _RAND_650;
  reg [31:0] mem_651;
  reg [31:0] _RAND_651;
  reg [31:0] mem_652;
  reg [31:0] _RAND_652;
  reg [31:0] mem_653;
  reg [31:0] _RAND_653;
  reg [31:0] mem_654;
  reg [31:0] _RAND_654;
  reg [31:0] mem_655;
  reg [31:0] _RAND_655;
  reg [31:0] mem_656;
  reg [31:0] _RAND_656;
  reg [31:0] mem_657;
  reg [31:0] _RAND_657;
  reg [31:0] mem_658;
  reg [31:0] _RAND_658;
  reg [31:0] mem_659;
  reg [31:0] _RAND_659;
  reg [31:0] mem_660;
  reg [31:0] _RAND_660;
  reg [31:0] mem_661;
  reg [31:0] _RAND_661;
  reg [31:0] mem_662;
  reg [31:0] _RAND_662;
  reg [31:0] mem_663;
  reg [31:0] _RAND_663;
  reg [31:0] mem_664;
  reg [31:0] _RAND_664;
  reg [31:0] mem_665;
  reg [31:0] _RAND_665;
  reg [31:0] mem_666;
  reg [31:0] _RAND_666;
  reg [31:0] mem_667;
  reg [31:0] _RAND_667;
  reg [31:0] mem_668;
  reg [31:0] _RAND_668;
  reg [31:0] mem_669;
  reg [31:0] _RAND_669;
  reg [31:0] mem_670;
  reg [31:0] _RAND_670;
  reg [31:0] mem_671;
  reg [31:0] _RAND_671;
  reg [31:0] mem_672;
  reg [31:0] _RAND_672;
  reg [31:0] mem_673;
  reg [31:0] _RAND_673;
  reg [31:0] mem_674;
  reg [31:0] _RAND_674;
  reg [31:0] mem_675;
  reg [31:0] _RAND_675;
  reg [31:0] mem_676;
  reg [31:0] _RAND_676;
  reg [31:0] mem_677;
  reg [31:0] _RAND_677;
  reg [31:0] mem_678;
  reg [31:0] _RAND_678;
  reg [31:0] mem_679;
  reg [31:0] _RAND_679;
  reg [31:0] mem_680;
  reg [31:0] _RAND_680;
  reg [31:0] mem_681;
  reg [31:0] _RAND_681;
  reg [31:0] mem_682;
  reg [31:0] _RAND_682;
  reg [31:0] mem_683;
  reg [31:0] _RAND_683;
  reg [31:0] mem_684;
  reg [31:0] _RAND_684;
  reg [31:0] mem_685;
  reg [31:0] _RAND_685;
  reg [31:0] mem_686;
  reg [31:0] _RAND_686;
  reg [31:0] mem_687;
  reg [31:0] _RAND_687;
  reg [31:0] mem_688;
  reg [31:0] _RAND_688;
  reg [31:0] mem_689;
  reg [31:0] _RAND_689;
  reg [31:0] mem_690;
  reg [31:0] _RAND_690;
  reg [31:0] mem_691;
  reg [31:0] _RAND_691;
  reg [31:0] mem_692;
  reg [31:0] _RAND_692;
  reg [31:0] mem_693;
  reg [31:0] _RAND_693;
  reg [31:0] mem_694;
  reg [31:0] _RAND_694;
  reg [31:0] mem_695;
  reg [31:0] _RAND_695;
  reg [31:0] mem_696;
  reg [31:0] _RAND_696;
  reg [31:0] mem_697;
  reg [31:0] _RAND_697;
  reg [31:0] mem_698;
  reg [31:0] _RAND_698;
  reg [31:0] mem_699;
  reg [31:0] _RAND_699;
  reg [31:0] mem_700;
  reg [31:0] _RAND_700;
  reg [31:0] mem_701;
  reg [31:0] _RAND_701;
  reg [31:0] mem_702;
  reg [31:0] _RAND_702;
  reg [31:0] mem_703;
  reg [31:0] _RAND_703;
  reg [31:0] mem_704;
  reg [31:0] _RAND_704;
  reg [31:0] mem_705;
  reg [31:0] _RAND_705;
  reg [31:0] mem_706;
  reg [31:0] _RAND_706;
  reg [31:0] mem_707;
  reg [31:0] _RAND_707;
  reg [31:0] mem_708;
  reg [31:0] _RAND_708;
  reg [31:0] mem_709;
  reg [31:0] _RAND_709;
  reg [31:0] mem_710;
  reg [31:0] _RAND_710;
  reg [31:0] mem_711;
  reg [31:0] _RAND_711;
  reg [31:0] mem_712;
  reg [31:0] _RAND_712;
  reg [31:0] mem_713;
  reg [31:0] _RAND_713;
  reg [31:0] mem_714;
  reg [31:0] _RAND_714;
  reg [31:0] mem_715;
  reg [31:0] _RAND_715;
  reg [31:0] mem_716;
  reg [31:0] _RAND_716;
  reg [31:0] mem_717;
  reg [31:0] _RAND_717;
  reg [31:0] mem_718;
  reg [31:0] _RAND_718;
  reg [31:0] mem_719;
  reg [31:0] _RAND_719;
  reg [31:0] mem_720;
  reg [31:0] _RAND_720;
  reg [31:0] mem_721;
  reg [31:0] _RAND_721;
  reg [31:0] mem_722;
  reg [31:0] _RAND_722;
  reg [31:0] mem_723;
  reg [31:0] _RAND_723;
  reg [31:0] mem_724;
  reg [31:0] _RAND_724;
  reg [31:0] mem_725;
  reg [31:0] _RAND_725;
  reg [31:0] mem_726;
  reg [31:0] _RAND_726;
  reg [31:0] mem_727;
  reg [31:0] _RAND_727;
  reg [31:0] mem_728;
  reg [31:0] _RAND_728;
  reg [31:0] mem_729;
  reg [31:0] _RAND_729;
  reg [31:0] mem_730;
  reg [31:0] _RAND_730;
  reg [31:0] mem_731;
  reg [31:0] _RAND_731;
  reg [31:0] mem_732;
  reg [31:0] _RAND_732;
  reg [31:0] mem_733;
  reg [31:0] _RAND_733;
  reg [31:0] mem_734;
  reg [31:0] _RAND_734;
  reg [31:0] mem_735;
  reg [31:0] _RAND_735;
  reg [31:0] mem_736;
  reg [31:0] _RAND_736;
  reg [31:0] mem_737;
  reg [31:0] _RAND_737;
  reg [31:0] mem_738;
  reg [31:0] _RAND_738;
  reg [31:0] mem_739;
  reg [31:0] _RAND_739;
  reg [31:0] mem_740;
  reg [31:0] _RAND_740;
  reg [31:0] mem_741;
  reg [31:0] _RAND_741;
  reg [31:0] mem_742;
  reg [31:0] _RAND_742;
  reg [31:0] mem_743;
  reg [31:0] _RAND_743;
  reg [31:0] mem_744;
  reg [31:0] _RAND_744;
  reg [31:0] mem_745;
  reg [31:0] _RAND_745;
  reg [31:0] mem_746;
  reg [31:0] _RAND_746;
  reg [31:0] mem_747;
  reg [31:0] _RAND_747;
  reg [31:0] mem_748;
  reg [31:0] _RAND_748;
  reg [31:0] mem_749;
  reg [31:0] _RAND_749;
  reg [31:0] mem_750;
  reg [31:0] _RAND_750;
  reg [31:0] mem_751;
  reg [31:0] _RAND_751;
  reg [31:0] mem_752;
  reg [31:0] _RAND_752;
  reg [31:0] mem_753;
  reg [31:0] _RAND_753;
  reg [31:0] mem_754;
  reg [31:0] _RAND_754;
  reg [31:0] mem_755;
  reg [31:0] _RAND_755;
  reg [31:0] mem_756;
  reg [31:0] _RAND_756;
  reg [31:0] mem_757;
  reg [31:0] _RAND_757;
  reg [31:0] mem_758;
  reg [31:0] _RAND_758;
  reg [31:0] mem_759;
  reg [31:0] _RAND_759;
  reg [31:0] mem_760;
  reg [31:0] _RAND_760;
  reg [31:0] mem_761;
  reg [31:0] _RAND_761;
  reg [31:0] mem_762;
  reg [31:0] _RAND_762;
  reg [31:0] mem_763;
  reg [31:0] _RAND_763;
  reg [31:0] mem_764;
  reg [31:0] _RAND_764;
  reg [31:0] mem_765;
  reg [31:0] _RAND_765;
  reg [31:0] mem_766;
  reg [31:0] _RAND_766;
  reg [31:0] mem_767;
  reg [31:0] _RAND_767;
  reg [31:0] mem_768;
  reg [31:0] _RAND_768;
  reg [31:0] mem_769;
  reg [31:0] _RAND_769;
  reg [31:0] mem_770;
  reg [31:0] _RAND_770;
  reg [31:0] mem_771;
  reg [31:0] _RAND_771;
  reg [31:0] mem_772;
  reg [31:0] _RAND_772;
  reg [31:0] mem_773;
  reg [31:0] _RAND_773;
  reg [31:0] mem_774;
  reg [31:0] _RAND_774;
  reg [31:0] mem_775;
  reg [31:0] _RAND_775;
  reg [31:0] mem_776;
  reg [31:0] _RAND_776;
  reg [31:0] mem_777;
  reg [31:0] _RAND_777;
  reg [31:0] mem_778;
  reg [31:0] _RAND_778;
  reg [31:0] mem_779;
  reg [31:0] _RAND_779;
  reg [31:0] mem_780;
  reg [31:0] _RAND_780;
  reg [31:0] mem_781;
  reg [31:0] _RAND_781;
  reg [31:0] mem_782;
  reg [31:0] _RAND_782;
  reg [31:0] mem_783;
  reg [31:0] _RAND_783;
  reg [31:0] mem_784;
  reg [31:0] _RAND_784;
  reg [31:0] mem_785;
  reg [31:0] _RAND_785;
  reg [31:0] mem_786;
  reg [31:0] _RAND_786;
  reg [31:0] mem_787;
  reg [31:0] _RAND_787;
  reg [31:0] mem_788;
  reg [31:0] _RAND_788;
  reg [31:0] mem_789;
  reg [31:0] _RAND_789;
  reg [31:0] mem_790;
  reg [31:0] _RAND_790;
  reg [31:0] mem_791;
  reg [31:0] _RAND_791;
  reg [31:0] mem_792;
  reg [31:0] _RAND_792;
  reg [31:0] mem_793;
  reg [31:0] _RAND_793;
  reg [31:0] mem_794;
  reg [31:0] _RAND_794;
  reg [31:0] mem_795;
  reg [31:0] _RAND_795;
  reg [31:0] mem_796;
  reg [31:0] _RAND_796;
  reg [31:0] mem_797;
  reg [31:0] _RAND_797;
  reg [31:0] mem_798;
  reg [31:0] _RAND_798;
  reg [31:0] mem_799;
  reg [31:0] _RAND_799;
  reg [31:0] mem_800;
  reg [31:0] _RAND_800;
  reg [31:0] mem_801;
  reg [31:0] _RAND_801;
  reg [31:0] mem_802;
  reg [31:0] _RAND_802;
  reg [31:0] mem_803;
  reg [31:0] _RAND_803;
  reg [31:0] mem_804;
  reg [31:0] _RAND_804;
  reg [31:0] mem_805;
  reg [31:0] _RAND_805;
  reg [31:0] mem_806;
  reg [31:0] _RAND_806;
  reg [31:0] mem_807;
  reg [31:0] _RAND_807;
  reg [31:0] mem_808;
  reg [31:0] _RAND_808;
  reg [31:0] mem_809;
  reg [31:0] _RAND_809;
  reg [31:0] mem_810;
  reg [31:0] _RAND_810;
  reg [31:0] mem_811;
  reg [31:0] _RAND_811;
  reg [31:0] mem_812;
  reg [31:0] _RAND_812;
  reg [31:0] mem_813;
  reg [31:0] _RAND_813;
  reg [31:0] mem_814;
  reg [31:0] _RAND_814;
  reg [31:0] mem_815;
  reg [31:0] _RAND_815;
  reg [31:0] mem_816;
  reg [31:0] _RAND_816;
  reg [31:0] mem_817;
  reg [31:0] _RAND_817;
  reg [31:0] mem_818;
  reg [31:0] _RAND_818;
  reg [31:0] mem_819;
  reg [31:0] _RAND_819;
  reg [31:0] mem_820;
  reg [31:0] _RAND_820;
  reg [31:0] mem_821;
  reg [31:0] _RAND_821;
  reg [31:0] mem_822;
  reg [31:0] _RAND_822;
  reg [31:0] mem_823;
  reg [31:0] _RAND_823;
  reg [31:0] mem_824;
  reg [31:0] _RAND_824;
  reg [31:0] mem_825;
  reg [31:0] _RAND_825;
  reg [31:0] mem_826;
  reg [31:0] _RAND_826;
  reg [31:0] mem_827;
  reg [31:0] _RAND_827;
  reg [31:0] mem_828;
  reg [31:0] _RAND_828;
  reg [31:0] mem_829;
  reg [31:0] _RAND_829;
  reg [31:0] mem_830;
  reg [31:0] _RAND_830;
  reg [31:0] mem_831;
  reg [31:0] _RAND_831;
  reg [31:0] mem_832;
  reg [31:0] _RAND_832;
  reg [31:0] mem_833;
  reg [31:0] _RAND_833;
  reg [31:0] mem_834;
  reg [31:0] _RAND_834;
  reg [31:0] mem_835;
  reg [31:0] _RAND_835;
  reg [31:0] mem_836;
  reg [31:0] _RAND_836;
  reg [31:0] mem_837;
  reg [31:0] _RAND_837;
  reg [31:0] mem_838;
  reg [31:0] _RAND_838;
  reg [31:0] mem_839;
  reg [31:0] _RAND_839;
  reg [31:0] mem_840;
  reg [31:0] _RAND_840;
  reg [31:0] mem_841;
  reg [31:0] _RAND_841;
  reg [31:0] mem_842;
  reg [31:0] _RAND_842;
  reg [31:0] mem_843;
  reg [31:0] _RAND_843;
  reg [31:0] mem_844;
  reg [31:0] _RAND_844;
  reg [31:0] mem_845;
  reg [31:0] _RAND_845;
  reg [31:0] mem_846;
  reg [31:0] _RAND_846;
  reg [31:0] mem_847;
  reg [31:0] _RAND_847;
  reg [31:0] mem_848;
  reg [31:0] _RAND_848;
  reg [31:0] mem_849;
  reg [31:0] _RAND_849;
  reg [31:0] mem_850;
  reg [31:0] _RAND_850;
  reg [31:0] mem_851;
  reg [31:0] _RAND_851;
  reg [31:0] mem_852;
  reg [31:0] _RAND_852;
  reg [31:0] mem_853;
  reg [31:0] _RAND_853;
  reg [31:0] mem_854;
  reg [31:0] _RAND_854;
  reg [31:0] mem_855;
  reg [31:0] _RAND_855;
  reg [31:0] mem_856;
  reg [31:0] _RAND_856;
  reg [31:0] mem_857;
  reg [31:0] _RAND_857;
  reg [31:0] mem_858;
  reg [31:0] _RAND_858;
  reg [31:0] mem_859;
  reg [31:0] _RAND_859;
  reg [31:0] mem_860;
  reg [31:0] _RAND_860;
  reg [31:0] mem_861;
  reg [31:0] _RAND_861;
  reg [31:0] mem_862;
  reg [31:0] _RAND_862;
  reg [31:0] mem_863;
  reg [31:0] _RAND_863;
  reg [31:0] mem_864;
  reg [31:0] _RAND_864;
  reg [31:0] mem_865;
  reg [31:0] _RAND_865;
  reg [31:0] mem_866;
  reg [31:0] _RAND_866;
  reg [31:0] mem_867;
  reg [31:0] _RAND_867;
  reg [31:0] mem_868;
  reg [31:0] _RAND_868;
  reg [31:0] mem_869;
  reg [31:0] _RAND_869;
  reg [31:0] mem_870;
  reg [31:0] _RAND_870;
  reg [31:0] mem_871;
  reg [31:0] _RAND_871;
  reg [31:0] mem_872;
  reg [31:0] _RAND_872;
  reg [31:0] mem_873;
  reg [31:0] _RAND_873;
  reg [31:0] mem_874;
  reg [31:0] _RAND_874;
  reg [31:0] mem_875;
  reg [31:0] _RAND_875;
  reg [31:0] mem_876;
  reg [31:0] _RAND_876;
  reg [31:0] mem_877;
  reg [31:0] _RAND_877;
  reg [31:0] mem_878;
  reg [31:0] _RAND_878;
  reg [31:0] mem_879;
  reg [31:0] _RAND_879;
  reg [31:0] mem_880;
  reg [31:0] _RAND_880;
  reg [31:0] mem_881;
  reg [31:0] _RAND_881;
  reg [31:0] mem_882;
  reg [31:0] _RAND_882;
  reg [31:0] mem_883;
  reg [31:0] _RAND_883;
  reg [31:0] mem_884;
  reg [31:0] _RAND_884;
  reg [31:0] mem_885;
  reg [31:0] _RAND_885;
  reg [31:0] mem_886;
  reg [31:0] _RAND_886;
  reg [31:0] mem_887;
  reg [31:0] _RAND_887;
  reg [31:0] mem_888;
  reg [31:0] _RAND_888;
  reg [31:0] mem_889;
  reg [31:0] _RAND_889;
  reg [31:0] mem_890;
  reg [31:0] _RAND_890;
  reg [31:0] mem_891;
  reg [31:0] _RAND_891;
  reg [31:0] mem_892;
  reg [31:0] _RAND_892;
  reg [31:0] mem_893;
  reg [31:0] _RAND_893;
  reg [31:0] mem_894;
  reg [31:0] _RAND_894;
  reg [31:0] mem_895;
  reg [31:0] _RAND_895;
  reg [31:0] mem_896;
  reg [31:0] _RAND_896;
  reg [31:0] mem_897;
  reg [31:0] _RAND_897;
  reg [31:0] mem_898;
  reg [31:0] _RAND_898;
  reg [31:0] mem_899;
  reg [31:0] _RAND_899;
  reg [31:0] mem_900;
  reg [31:0] _RAND_900;
  reg [31:0] mem_901;
  reg [31:0] _RAND_901;
  reg [31:0] mem_902;
  reg [31:0] _RAND_902;
  reg [31:0] mem_903;
  reg [31:0] _RAND_903;
  reg [31:0] mem_904;
  reg [31:0] _RAND_904;
  reg [31:0] mem_905;
  reg [31:0] _RAND_905;
  reg [31:0] mem_906;
  reg [31:0] _RAND_906;
  reg [31:0] mem_907;
  reg [31:0] _RAND_907;
  reg [31:0] mem_908;
  reg [31:0] _RAND_908;
  reg [31:0] mem_909;
  reg [31:0] _RAND_909;
  reg [31:0] mem_910;
  reg [31:0] _RAND_910;
  reg [31:0] mem_911;
  reg [31:0] _RAND_911;
  reg [31:0] mem_912;
  reg [31:0] _RAND_912;
  reg [31:0] mem_913;
  reg [31:0] _RAND_913;
  reg [31:0] mem_914;
  reg [31:0] _RAND_914;
  reg [31:0] mem_915;
  reg [31:0] _RAND_915;
  reg [31:0] mem_916;
  reg [31:0] _RAND_916;
  reg [31:0] mem_917;
  reg [31:0] _RAND_917;
  reg [31:0] mem_918;
  reg [31:0] _RAND_918;
  reg [31:0] mem_919;
  reg [31:0] _RAND_919;
  reg [31:0] mem_920;
  reg [31:0] _RAND_920;
  reg [31:0] mem_921;
  reg [31:0] _RAND_921;
  reg [31:0] mem_922;
  reg [31:0] _RAND_922;
  reg [31:0] mem_923;
  reg [31:0] _RAND_923;
  reg [31:0] mem_924;
  reg [31:0] _RAND_924;
  reg [31:0] mem_925;
  reg [31:0] _RAND_925;
  reg [31:0] mem_926;
  reg [31:0] _RAND_926;
  reg [31:0] mem_927;
  reg [31:0] _RAND_927;
  reg [31:0] mem_928;
  reg [31:0] _RAND_928;
  reg [31:0] mem_929;
  reg [31:0] _RAND_929;
  reg [31:0] mem_930;
  reg [31:0] _RAND_930;
  reg [31:0] mem_931;
  reg [31:0] _RAND_931;
  reg [31:0] mem_932;
  reg [31:0] _RAND_932;
  reg [31:0] mem_933;
  reg [31:0] _RAND_933;
  reg [31:0] mem_934;
  reg [31:0] _RAND_934;
  reg [31:0] mem_935;
  reg [31:0] _RAND_935;
  reg [31:0] mem_936;
  reg [31:0] _RAND_936;
  reg [31:0] mem_937;
  reg [31:0] _RAND_937;
  reg [31:0] mem_938;
  reg [31:0] _RAND_938;
  reg [31:0] mem_939;
  reg [31:0] _RAND_939;
  reg [31:0] mem_940;
  reg [31:0] _RAND_940;
  reg [31:0] mem_941;
  reg [31:0] _RAND_941;
  reg [31:0] mem_942;
  reg [31:0] _RAND_942;
  reg [31:0] mem_943;
  reg [31:0] _RAND_943;
  reg [31:0] mem_944;
  reg [31:0] _RAND_944;
  reg [31:0] mem_945;
  reg [31:0] _RAND_945;
  reg [31:0] mem_946;
  reg [31:0] _RAND_946;
  reg [31:0] mem_947;
  reg [31:0] _RAND_947;
  reg [31:0] mem_948;
  reg [31:0] _RAND_948;
  reg [31:0] mem_949;
  reg [31:0] _RAND_949;
  reg [31:0] mem_950;
  reg [31:0] _RAND_950;
  reg [31:0] mem_951;
  reg [31:0] _RAND_951;
  reg [31:0] mem_952;
  reg [31:0] _RAND_952;
  reg [31:0] mem_953;
  reg [31:0] _RAND_953;
  reg [31:0] mem_954;
  reg [31:0] _RAND_954;
  reg [31:0] mem_955;
  reg [31:0] _RAND_955;
  reg [31:0] mem_956;
  reg [31:0] _RAND_956;
  reg [31:0] mem_957;
  reg [31:0] _RAND_957;
  reg [31:0] mem_958;
  reg [31:0] _RAND_958;
  reg [31:0] mem_959;
  reg [31:0] _RAND_959;
  reg [31:0] mem_960;
  reg [31:0] _RAND_960;
  reg [31:0] mem_961;
  reg [31:0] _RAND_961;
  reg [31:0] mem_962;
  reg [31:0] _RAND_962;
  reg [31:0] mem_963;
  reg [31:0] _RAND_963;
  reg [31:0] mem_964;
  reg [31:0] _RAND_964;
  reg [31:0] mem_965;
  reg [31:0] _RAND_965;
  reg [31:0] mem_966;
  reg [31:0] _RAND_966;
  reg [31:0] mem_967;
  reg [31:0] _RAND_967;
  reg [31:0] mem_968;
  reg [31:0] _RAND_968;
  reg [31:0] mem_969;
  reg [31:0] _RAND_969;
  reg [31:0] mem_970;
  reg [31:0] _RAND_970;
  reg [31:0] mem_971;
  reg [31:0] _RAND_971;
  reg [31:0] mem_972;
  reg [31:0] _RAND_972;
  reg [31:0] mem_973;
  reg [31:0] _RAND_973;
  reg [31:0] mem_974;
  reg [31:0] _RAND_974;
  reg [31:0] mem_975;
  reg [31:0] _RAND_975;
  reg [31:0] mem_976;
  reg [31:0] _RAND_976;
  reg [31:0] mem_977;
  reg [31:0] _RAND_977;
  reg [31:0] mem_978;
  reg [31:0] _RAND_978;
  reg [31:0] mem_979;
  reg [31:0] _RAND_979;
  reg [31:0] mem_980;
  reg [31:0] _RAND_980;
  reg [31:0] mem_981;
  reg [31:0] _RAND_981;
  reg [31:0] mem_982;
  reg [31:0] _RAND_982;
  reg [31:0] mem_983;
  reg [31:0] _RAND_983;
  reg [31:0] mem_984;
  reg [31:0] _RAND_984;
  reg [31:0] mem_985;
  reg [31:0] _RAND_985;
  reg [31:0] mem_986;
  reg [31:0] _RAND_986;
  reg [31:0] mem_987;
  reg [31:0] _RAND_987;
  reg [31:0] mem_988;
  reg [31:0] _RAND_988;
  reg [31:0] mem_989;
  reg [31:0] _RAND_989;
  reg [31:0] mem_990;
  reg [31:0] _RAND_990;
  reg [31:0] mem_991;
  reg [31:0] _RAND_991;
  reg [31:0] mem_992;
  reg [31:0] _RAND_992;
  reg [31:0] mem_993;
  reg [31:0] _RAND_993;
  reg [31:0] mem_994;
  reg [31:0] _RAND_994;
  reg [31:0] mem_995;
  reg [31:0] _RAND_995;
  reg [31:0] mem_996;
  reg [31:0] _RAND_996;
  reg [31:0] mem_997;
  reg [31:0] _RAND_997;
  reg [31:0] mem_998;
  reg [31:0] _RAND_998;
  reg [31:0] mem_999;
  reg [31:0] _RAND_999;
  reg [31:0] mem_1000;
  reg [31:0] _RAND_1000;
  reg [31:0] mem_1001;
  reg [31:0] _RAND_1001;
  reg [31:0] mem_1002;
  reg [31:0] _RAND_1002;
  reg [31:0] mem_1003;
  reg [31:0] _RAND_1003;
  reg [31:0] mem_1004;
  reg [31:0] _RAND_1004;
  reg [31:0] mem_1005;
  reg [31:0] _RAND_1005;
  reg [31:0] mem_1006;
  reg [31:0] _RAND_1006;
  reg [31:0] mem_1007;
  reg [31:0] _RAND_1007;
  reg [31:0] mem_1008;
  reg [31:0] _RAND_1008;
  reg [31:0] mem_1009;
  reg [31:0] _RAND_1009;
  reg [31:0] mem_1010;
  reg [31:0] _RAND_1010;
  reg [31:0] mem_1011;
  reg [31:0] _RAND_1011;
  reg [31:0] mem_1012;
  reg [31:0] _RAND_1012;
  reg [31:0] mem_1013;
  reg [31:0] _RAND_1013;
  reg [31:0] mem_1014;
  reg [31:0] _RAND_1014;
  reg [31:0] mem_1015;
  reg [31:0] _RAND_1015;
  reg [31:0] mem_1016;
  reg [31:0] _RAND_1016;
  reg [31:0] mem_1017;
  reg [31:0] _RAND_1017;
  reg [31:0] mem_1018;
  reg [31:0] _RAND_1018;
  reg [31:0] mem_1019;
  reg [31:0] _RAND_1019;
  reg [31:0] mem_1020;
  reg [31:0] _RAND_1020;
  reg [31:0] mem_1021;
  reg [31:0] _RAND_1021;
  reg [31:0] mem_1022;
  reg [31:0] _RAND_1022;
  reg [31:0] mem_1023;
  reg [31:0] _RAND_1023;
  reg [31:0] mem_1024;
  reg [31:0] _RAND_1024;
  reg [31:0] mem_1025;
  reg [31:0] _RAND_1025;
  reg [31:0] mem_1026;
  reg [31:0] _RAND_1026;
  reg [31:0] mem_1027;
  reg [31:0] _RAND_1027;
  reg [31:0] mem_1028;
  reg [31:0] _RAND_1028;
  reg [31:0] mem_1029;
  reg [31:0] _RAND_1029;
  reg [31:0] mem_1030;
  reg [31:0] _RAND_1030;
  reg [31:0] mem_1031;
  reg [31:0] _RAND_1031;
  reg [31:0] mem_1032;
  reg [31:0] _RAND_1032;
  reg [31:0] mem_1033;
  reg [31:0] _RAND_1033;
  reg [31:0] mem_1034;
  reg [31:0] _RAND_1034;
  reg [31:0] mem_1035;
  reg [31:0] _RAND_1035;
  reg [31:0] mem_1036;
  reg [31:0] _RAND_1036;
  reg [31:0] mem_1037;
  reg [31:0] _RAND_1037;
  reg [31:0] mem_1038;
  reg [31:0] _RAND_1038;
  reg [31:0] mem_1039;
  reg [31:0] _RAND_1039;
  reg [31:0] mem_1040;
  reg [31:0] _RAND_1040;
  reg [31:0] mem_1041;
  reg [31:0] _RAND_1041;
  reg [31:0] mem_1042;
  reg [31:0] _RAND_1042;
  reg [31:0] mem_1043;
  reg [31:0] _RAND_1043;
  reg [31:0] mem_1044;
  reg [31:0] _RAND_1044;
  reg [31:0] mem_1045;
  reg [31:0] _RAND_1045;
  reg [31:0] mem_1046;
  reg [31:0] _RAND_1046;
  reg [31:0] mem_1047;
  reg [31:0] _RAND_1047;
  reg [31:0] mem_1048;
  reg [31:0] _RAND_1048;
  reg [31:0] mem_1049;
  reg [31:0] _RAND_1049;
  reg [31:0] mem_1050;
  reg [31:0] _RAND_1050;
  reg [31:0] mem_1051;
  reg [31:0] _RAND_1051;
  reg [31:0] mem_1052;
  reg [31:0] _RAND_1052;
  reg [31:0] mem_1053;
  reg [31:0] _RAND_1053;
  reg [31:0] mem_1054;
  reg [31:0] _RAND_1054;
  reg [31:0] mem_1055;
  reg [31:0] _RAND_1055;
  reg [31:0] mem_1056;
  reg [31:0] _RAND_1056;
  reg [31:0] mem_1057;
  reg [31:0] _RAND_1057;
  reg [31:0] mem_1058;
  reg [31:0] _RAND_1058;
  reg [31:0] mem_1059;
  reg [31:0] _RAND_1059;
  reg [31:0] mem_1060;
  reg [31:0] _RAND_1060;
  reg [31:0] mem_1061;
  reg [31:0] _RAND_1061;
  reg [31:0] mem_1062;
  reg [31:0] _RAND_1062;
  reg [31:0] mem_1063;
  reg [31:0] _RAND_1063;
  reg [31:0] mem_1064;
  reg [31:0] _RAND_1064;
  reg [31:0] mem_1065;
  reg [31:0] _RAND_1065;
  reg [31:0] mem_1066;
  reg [31:0] _RAND_1066;
  reg [31:0] mem_1067;
  reg [31:0] _RAND_1067;
  reg [31:0] mem_1068;
  reg [31:0] _RAND_1068;
  reg [31:0] mem_1069;
  reg [31:0] _RAND_1069;
  reg [31:0] mem_1070;
  reg [31:0] _RAND_1070;
  reg [31:0] mem_1071;
  reg [31:0] _RAND_1071;
  reg [31:0] mem_1072;
  reg [31:0] _RAND_1072;
  reg [31:0] mem_1073;
  reg [31:0] _RAND_1073;
  reg [31:0] mem_1074;
  reg [31:0] _RAND_1074;
  reg [31:0] mem_1075;
  reg [31:0] _RAND_1075;
  reg [31:0] mem_1076;
  reg [31:0] _RAND_1076;
  reg [31:0] mem_1077;
  reg [31:0] _RAND_1077;
  reg [31:0] mem_1078;
  reg [31:0] _RAND_1078;
  reg [31:0] mem_1079;
  reg [31:0] _RAND_1079;
  reg [31:0] mem_1080;
  reg [31:0] _RAND_1080;
  reg [31:0] mem_1081;
  reg [31:0] _RAND_1081;
  reg [31:0] mem_1082;
  reg [31:0] _RAND_1082;
  reg [31:0] mem_1083;
  reg [31:0] _RAND_1083;
  reg [31:0] mem_1084;
  reg [31:0] _RAND_1084;
  reg [31:0] mem_1085;
  reg [31:0] _RAND_1085;
  reg [31:0] mem_1086;
  reg [31:0] _RAND_1086;
  reg [31:0] mem_1087;
  reg [31:0] _RAND_1087;
  reg [31:0] mem_1088;
  reg [31:0] _RAND_1088;
  reg [31:0] mem_1089;
  reg [31:0] _RAND_1089;
  reg [31:0] mem_1090;
  reg [31:0] _RAND_1090;
  reg [31:0] mem_1091;
  reg [31:0] _RAND_1091;
  reg [31:0] mem_1092;
  reg [31:0] _RAND_1092;
  reg [31:0] mem_1093;
  reg [31:0] _RAND_1093;
  reg [31:0] mem_1094;
  reg [31:0] _RAND_1094;
  reg [31:0] mem_1095;
  reg [31:0] _RAND_1095;
  reg [31:0] mem_1096;
  reg [31:0] _RAND_1096;
  reg [31:0] mem_1097;
  reg [31:0] _RAND_1097;
  reg [31:0] mem_1098;
  reg [31:0] _RAND_1098;
  reg [31:0] mem_1099;
  reg [31:0] _RAND_1099;
  reg [31:0] mem_1100;
  reg [31:0] _RAND_1100;
  reg [31:0] mem_1101;
  reg [31:0] _RAND_1101;
  reg [31:0] mem_1102;
  reg [31:0] _RAND_1102;
  reg [31:0] mem_1103;
  reg [31:0] _RAND_1103;
  reg [31:0] mem_1104;
  reg [31:0] _RAND_1104;
  reg [31:0] mem_1105;
  reg [31:0] _RAND_1105;
  reg [31:0] mem_1106;
  reg [31:0] _RAND_1106;
  reg [31:0] mem_1107;
  reg [31:0] _RAND_1107;
  reg [31:0] mem_1108;
  reg [31:0] _RAND_1108;
  reg [31:0] mem_1109;
  reg [31:0] _RAND_1109;
  reg [31:0] mem_1110;
  reg [31:0] _RAND_1110;
  reg [31:0] mem_1111;
  reg [31:0] _RAND_1111;
  reg [31:0] mem_1112;
  reg [31:0] _RAND_1112;
  reg [31:0] mem_1113;
  reg [31:0] _RAND_1113;
  reg [31:0] mem_1114;
  reg [31:0] _RAND_1114;
  reg [31:0] mem_1115;
  reg [31:0] _RAND_1115;
  reg [31:0] mem_1116;
  reg [31:0] _RAND_1116;
  reg [31:0] mem_1117;
  reg [31:0] _RAND_1117;
  reg [31:0] mem_1118;
  reg [31:0] _RAND_1118;
  reg [31:0] mem_1119;
  reg [31:0] _RAND_1119;
  reg [31:0] mem_1120;
  reg [31:0] _RAND_1120;
  reg [31:0] mem_1121;
  reg [31:0] _RAND_1121;
  reg [31:0] mem_1122;
  reg [31:0] _RAND_1122;
  reg [31:0] mem_1123;
  reg [31:0] _RAND_1123;
  reg [31:0] mem_1124;
  reg [31:0] _RAND_1124;
  reg [31:0] mem_1125;
  reg [31:0] _RAND_1125;
  reg [31:0] mem_1126;
  reg [31:0] _RAND_1126;
  reg [31:0] mem_1127;
  reg [31:0] _RAND_1127;
  reg [31:0] mem_1128;
  reg [31:0] _RAND_1128;
  reg [31:0] mem_1129;
  reg [31:0] _RAND_1129;
  reg [31:0] mem_1130;
  reg [31:0] _RAND_1130;
  reg [31:0] mem_1131;
  reg [31:0] _RAND_1131;
  reg [31:0] mem_1132;
  reg [31:0] _RAND_1132;
  reg [31:0] mem_1133;
  reg [31:0] _RAND_1133;
  reg [31:0] mem_1134;
  reg [31:0] _RAND_1134;
  reg [31:0] mem_1135;
  reg [31:0] _RAND_1135;
  reg [31:0] mem_1136;
  reg [31:0] _RAND_1136;
  reg [31:0] mem_1137;
  reg [31:0] _RAND_1137;
  reg [31:0] mem_1138;
  reg [31:0] _RAND_1138;
  reg [31:0] mem_1139;
  reg [31:0] _RAND_1139;
  reg [31:0] mem_1140;
  reg [31:0] _RAND_1140;
  reg [31:0] mem_1141;
  reg [31:0] _RAND_1141;
  reg [31:0] mem_1142;
  reg [31:0] _RAND_1142;
  reg [31:0] mem_1143;
  reg [31:0] _RAND_1143;
  reg [31:0] mem_1144;
  reg [31:0] _RAND_1144;
  reg [31:0] mem_1145;
  reg [31:0] _RAND_1145;
  reg [31:0] mem_1146;
  reg [31:0] _RAND_1146;
  reg [31:0] mem_1147;
  reg [31:0] _RAND_1147;
  reg [31:0] mem_1148;
  reg [31:0] _RAND_1148;
  reg [31:0] mem_1149;
  reg [31:0] _RAND_1149;
  reg [31:0] mem_1150;
  reg [31:0] _RAND_1150;
  reg [31:0] mem_1151;
  reg [31:0] _RAND_1151;
  reg [31:0] mem_1152;
  reg [31:0] _RAND_1152;
  reg [31:0] mem_1153;
  reg [31:0] _RAND_1153;
  reg [31:0] mem_1154;
  reg [31:0] _RAND_1154;
  reg [31:0] mem_1155;
  reg [31:0] _RAND_1155;
  reg [31:0] mem_1156;
  reg [31:0] _RAND_1156;
  reg [31:0] mem_1157;
  reg [31:0] _RAND_1157;
  reg [31:0] mem_1158;
  reg [31:0] _RAND_1158;
  reg [31:0] mem_1159;
  reg [31:0] _RAND_1159;
  reg [31:0] mem_1160;
  reg [31:0] _RAND_1160;
  reg [31:0] mem_1161;
  reg [31:0] _RAND_1161;
  reg [31:0] mem_1162;
  reg [31:0] _RAND_1162;
  reg [31:0] mem_1163;
  reg [31:0] _RAND_1163;
  reg [31:0] mem_1164;
  reg [31:0] _RAND_1164;
  reg [31:0] mem_1165;
  reg [31:0] _RAND_1165;
  reg [31:0] mem_1166;
  reg [31:0] _RAND_1166;
  reg [31:0] mem_1167;
  reg [31:0] _RAND_1167;
  reg [31:0] mem_1168;
  reg [31:0] _RAND_1168;
  reg [31:0] mem_1169;
  reg [31:0] _RAND_1169;
  reg [31:0] mem_1170;
  reg [31:0] _RAND_1170;
  reg [31:0] mem_1171;
  reg [31:0] _RAND_1171;
  reg [31:0] mem_1172;
  reg [31:0] _RAND_1172;
  reg [31:0] mem_1173;
  reg [31:0] _RAND_1173;
  reg [31:0] mem_1174;
  reg [31:0] _RAND_1174;
  reg [31:0] mem_1175;
  reg [31:0] _RAND_1175;
  reg [31:0] mem_1176;
  reg [31:0] _RAND_1176;
  reg [31:0] mem_1177;
  reg [31:0] _RAND_1177;
  reg [31:0] mem_1178;
  reg [31:0] _RAND_1178;
  reg [31:0] mem_1179;
  reg [31:0] _RAND_1179;
  reg [31:0] mem_1180;
  reg [31:0] _RAND_1180;
  reg [31:0] mem_1181;
  reg [31:0] _RAND_1181;
  reg [31:0] mem_1182;
  reg [31:0] _RAND_1182;
  reg [31:0] mem_1183;
  reg [31:0] _RAND_1183;
  reg [31:0] mem_1184;
  reg [31:0] _RAND_1184;
  reg [31:0] mem_1185;
  reg [31:0] _RAND_1185;
  reg [31:0] mem_1186;
  reg [31:0] _RAND_1186;
  reg [31:0] mem_1187;
  reg [31:0] _RAND_1187;
  reg [31:0] mem_1188;
  reg [31:0] _RAND_1188;
  reg [31:0] mem_1189;
  reg [31:0] _RAND_1189;
  reg [31:0] mem_1190;
  reg [31:0] _RAND_1190;
  reg [31:0] mem_1191;
  reg [31:0] _RAND_1191;
  reg [31:0] mem_1192;
  reg [31:0] _RAND_1192;
  reg [31:0] mem_1193;
  reg [31:0] _RAND_1193;
  reg [31:0] mem_1194;
  reg [31:0] _RAND_1194;
  reg [31:0] mem_1195;
  reg [31:0] _RAND_1195;
  reg [31:0] mem_1196;
  reg [31:0] _RAND_1196;
  reg [31:0] mem_1197;
  reg [31:0] _RAND_1197;
  reg [31:0] mem_1198;
  reg [31:0] _RAND_1198;
  reg [31:0] mem_1199;
  reg [31:0] _RAND_1199;
  reg [31:0] mem_1200;
  reg [31:0] _RAND_1200;
  reg [31:0] mem_1201;
  reg [31:0] _RAND_1201;
  reg [31:0] mem_1202;
  reg [31:0] _RAND_1202;
  reg [31:0] mem_1203;
  reg [31:0] _RAND_1203;
  reg [31:0] mem_1204;
  reg [31:0] _RAND_1204;
  reg [31:0] mem_1205;
  reg [31:0] _RAND_1205;
  reg [31:0] mem_1206;
  reg [31:0] _RAND_1206;
  reg [31:0] mem_1207;
  reg [31:0] _RAND_1207;
  reg [31:0] mem_1208;
  reg [31:0] _RAND_1208;
  reg [31:0] mem_1209;
  reg [31:0] _RAND_1209;
  reg [31:0] mem_1210;
  reg [31:0] _RAND_1210;
  reg [31:0] mem_1211;
  reg [31:0] _RAND_1211;
  reg [31:0] mem_1212;
  reg [31:0] _RAND_1212;
  reg [31:0] mem_1213;
  reg [31:0] _RAND_1213;
  reg [31:0] mem_1214;
  reg [31:0] _RAND_1214;
  reg [31:0] mem_1215;
  reg [31:0] _RAND_1215;
  reg [31:0] mem_1216;
  reg [31:0] _RAND_1216;
  reg [31:0] mem_1217;
  reg [31:0] _RAND_1217;
  reg [31:0] mem_1218;
  reg [31:0] _RAND_1218;
  reg [31:0] mem_1219;
  reg [31:0] _RAND_1219;
  reg [31:0] mem_1220;
  reg [31:0] _RAND_1220;
  reg [31:0] mem_1221;
  reg [31:0] _RAND_1221;
  reg [31:0] mem_1222;
  reg [31:0] _RAND_1222;
  reg [31:0] mem_1223;
  reg [31:0] _RAND_1223;
  reg [31:0] mem_1224;
  reg [31:0] _RAND_1224;
  reg [31:0] mem_1225;
  reg [31:0] _RAND_1225;
  reg [31:0] mem_1226;
  reg [31:0] _RAND_1226;
  reg [31:0] mem_1227;
  reg [31:0] _RAND_1227;
  reg [31:0] mem_1228;
  reg [31:0] _RAND_1228;
  reg [31:0] mem_1229;
  reg [31:0] _RAND_1229;
  reg [31:0] mem_1230;
  reg [31:0] _RAND_1230;
  reg [31:0] mem_1231;
  reg [31:0] _RAND_1231;
  reg [31:0] mem_1232;
  reg [31:0] _RAND_1232;
  reg [31:0] mem_1233;
  reg [31:0] _RAND_1233;
  reg [31:0] mem_1234;
  reg [31:0] _RAND_1234;
  reg [31:0] mem_1235;
  reg [31:0] _RAND_1235;
  reg [31:0] mem_1236;
  reg [31:0] _RAND_1236;
  reg [31:0] mem_1237;
  reg [31:0] _RAND_1237;
  reg [31:0] mem_1238;
  reg [31:0] _RAND_1238;
  reg [31:0] mem_1239;
  reg [31:0] _RAND_1239;
  reg [31:0] mem_1240;
  reg [31:0] _RAND_1240;
  reg [31:0] mem_1241;
  reg [31:0] _RAND_1241;
  reg [31:0] mem_1242;
  reg [31:0] _RAND_1242;
  reg [31:0] mem_1243;
  reg [31:0] _RAND_1243;
  reg [31:0] mem_1244;
  reg [31:0] _RAND_1244;
  reg [31:0] mem_1245;
  reg [31:0] _RAND_1245;
  reg [31:0] mem_1246;
  reg [31:0] _RAND_1246;
  reg [31:0] mem_1247;
  reg [31:0] _RAND_1247;
  reg [31:0] mem_1248;
  reg [31:0] _RAND_1248;
  reg [31:0] mem_1249;
  reg [31:0] _RAND_1249;
  reg [31:0] mem_1250;
  reg [31:0] _RAND_1250;
  reg [31:0] mem_1251;
  reg [31:0] _RAND_1251;
  reg [31:0] mem_1252;
  reg [31:0] _RAND_1252;
  reg [31:0] mem_1253;
  reg [31:0] _RAND_1253;
  reg [31:0] mem_1254;
  reg [31:0] _RAND_1254;
  reg [31:0] mem_1255;
  reg [31:0] _RAND_1255;
  reg [31:0] mem_1256;
  reg [31:0] _RAND_1256;
  reg [31:0] mem_1257;
  reg [31:0] _RAND_1257;
  reg [31:0] mem_1258;
  reg [31:0] _RAND_1258;
  reg [31:0] mem_1259;
  reg [31:0] _RAND_1259;
  reg [31:0] mem_1260;
  reg [31:0] _RAND_1260;
  reg [31:0] mem_1261;
  reg [31:0] _RAND_1261;
  reg [31:0] mem_1262;
  reg [31:0] _RAND_1262;
  reg [31:0] mem_1263;
  reg [31:0] _RAND_1263;
  reg [31:0] mem_1264;
  reg [31:0] _RAND_1264;
  reg [31:0] mem_1265;
  reg [31:0] _RAND_1265;
  reg [31:0] mem_1266;
  reg [31:0] _RAND_1266;
  reg [31:0] mem_1267;
  reg [31:0] _RAND_1267;
  reg [31:0] mem_1268;
  reg [31:0] _RAND_1268;
  reg [31:0] mem_1269;
  reg [31:0] _RAND_1269;
  reg [31:0] mem_1270;
  reg [31:0] _RAND_1270;
  reg [31:0] mem_1271;
  reg [31:0] _RAND_1271;
  reg [31:0] mem_1272;
  reg [31:0] _RAND_1272;
  reg [31:0] mem_1273;
  reg [31:0] _RAND_1273;
  reg [31:0] mem_1274;
  reg [31:0] _RAND_1274;
  reg [31:0] mem_1275;
  reg [31:0] _RAND_1275;
  reg [31:0] mem_1276;
  reg [31:0] _RAND_1276;
  reg [31:0] mem_1277;
  reg [31:0] _RAND_1277;
  reg [31:0] mem_1278;
  reg [31:0] _RAND_1278;
  reg [31:0] mem_1279;
  reg [31:0] _RAND_1279;
  reg [31:0] mem_1280;
  reg [31:0] _RAND_1280;
  reg [31:0] mem_1281;
  reg [31:0] _RAND_1281;
  reg [31:0] mem_1282;
  reg [31:0] _RAND_1282;
  reg [31:0] mem_1283;
  reg [31:0] _RAND_1283;
  reg [31:0] mem_1284;
  reg [31:0] _RAND_1284;
  reg [31:0] mem_1285;
  reg [31:0] _RAND_1285;
  reg [31:0] mem_1286;
  reg [31:0] _RAND_1286;
  reg [31:0] mem_1287;
  reg [31:0] _RAND_1287;
  reg [31:0] mem_1288;
  reg [31:0] _RAND_1288;
  reg [31:0] mem_1289;
  reg [31:0] _RAND_1289;
  reg [31:0] mem_1290;
  reg [31:0] _RAND_1290;
  reg [31:0] mem_1291;
  reg [31:0] _RAND_1291;
  reg [31:0] mem_1292;
  reg [31:0] _RAND_1292;
  reg [31:0] mem_1293;
  reg [31:0] _RAND_1293;
  reg [31:0] mem_1294;
  reg [31:0] _RAND_1294;
  reg [31:0] mem_1295;
  reg [31:0] _RAND_1295;
  reg [31:0] mem_1296;
  reg [31:0] _RAND_1296;
  reg [31:0] mem_1297;
  reg [31:0] _RAND_1297;
  reg [31:0] mem_1298;
  reg [31:0] _RAND_1298;
  reg [31:0] mem_1299;
  reg [31:0] _RAND_1299;
  reg [31:0] mem_1300;
  reg [31:0] _RAND_1300;
  reg [31:0] mem_1301;
  reg [31:0] _RAND_1301;
  reg [31:0] mem_1302;
  reg [31:0] _RAND_1302;
  reg [31:0] mem_1303;
  reg [31:0] _RAND_1303;
  reg [31:0] mem_1304;
  reg [31:0] _RAND_1304;
  reg [31:0] mem_1305;
  reg [31:0] _RAND_1305;
  reg [31:0] mem_1306;
  reg [31:0] _RAND_1306;
  reg [31:0] mem_1307;
  reg [31:0] _RAND_1307;
  reg [31:0] mem_1308;
  reg [31:0] _RAND_1308;
  reg [31:0] mem_1309;
  reg [31:0] _RAND_1309;
  reg [31:0] mem_1310;
  reg [31:0] _RAND_1310;
  reg [31:0] mem_1311;
  reg [31:0] _RAND_1311;
  reg [31:0] mem_1312;
  reg [31:0] _RAND_1312;
  reg [31:0] mem_1313;
  reg [31:0] _RAND_1313;
  reg [31:0] mem_1314;
  reg [31:0] _RAND_1314;
  reg [31:0] mem_1315;
  reg [31:0] _RAND_1315;
  reg [31:0] mem_1316;
  reg [31:0] _RAND_1316;
  reg [31:0] mem_1317;
  reg [31:0] _RAND_1317;
  reg [31:0] mem_1318;
  reg [31:0] _RAND_1318;
  reg [31:0] mem_1319;
  reg [31:0] _RAND_1319;
  reg [31:0] mem_1320;
  reg [31:0] _RAND_1320;
  reg [31:0] mem_1321;
  reg [31:0] _RAND_1321;
  reg [31:0] mem_1322;
  reg [31:0] _RAND_1322;
  reg [31:0] mem_1323;
  reg [31:0] _RAND_1323;
  reg [31:0] mem_1324;
  reg [31:0] _RAND_1324;
  reg [31:0] mem_1325;
  reg [31:0] _RAND_1325;
  reg [31:0] mem_1326;
  reg [31:0] _RAND_1326;
  reg [31:0] mem_1327;
  reg [31:0] _RAND_1327;
  reg [31:0] mem_1328;
  reg [31:0] _RAND_1328;
  reg [31:0] mem_1329;
  reg [31:0] _RAND_1329;
  reg [31:0] mem_1330;
  reg [31:0] _RAND_1330;
  reg [31:0] mem_1331;
  reg [31:0] _RAND_1331;
  reg [31:0] mem_1332;
  reg [31:0] _RAND_1332;
  reg [31:0] mem_1333;
  reg [31:0] _RAND_1333;
  reg [31:0] mem_1334;
  reg [31:0] _RAND_1334;
  reg [31:0] mem_1335;
  reg [31:0] _RAND_1335;
  reg [31:0] mem_1336;
  reg [31:0] _RAND_1336;
  reg [31:0] mem_1337;
  reg [31:0] _RAND_1337;
  reg [31:0] mem_1338;
  reg [31:0] _RAND_1338;
  reg [31:0] mem_1339;
  reg [31:0] _RAND_1339;
  reg [31:0] mem_1340;
  reg [31:0] _RAND_1340;
  reg [31:0] mem_1341;
  reg [31:0] _RAND_1341;
  reg [31:0] mem_1342;
  reg [31:0] _RAND_1342;
  reg [31:0] mem_1343;
  reg [31:0] _RAND_1343;
  reg [31:0] mem_1344;
  reg [31:0] _RAND_1344;
  reg [31:0] mem_1345;
  reg [31:0] _RAND_1345;
  reg [31:0] mem_1346;
  reg [31:0] _RAND_1346;
  reg [31:0] mem_1347;
  reg [31:0] _RAND_1347;
  reg [31:0] mem_1348;
  reg [31:0] _RAND_1348;
  reg [31:0] mem_1349;
  reg [31:0] _RAND_1349;
  reg [31:0] mem_1350;
  reg [31:0] _RAND_1350;
  reg [31:0] mem_1351;
  reg [31:0] _RAND_1351;
  reg [31:0] mem_1352;
  reg [31:0] _RAND_1352;
  reg [31:0] mem_1353;
  reg [31:0] _RAND_1353;
  reg [31:0] mem_1354;
  reg [31:0] _RAND_1354;
  reg [31:0] mem_1355;
  reg [31:0] _RAND_1355;
  reg [31:0] mem_1356;
  reg [31:0] _RAND_1356;
  reg [31:0] mem_1357;
  reg [31:0] _RAND_1357;
  reg [31:0] mem_1358;
  reg [31:0] _RAND_1358;
  reg [31:0] mem_1359;
  reg [31:0] _RAND_1359;
  reg [31:0] mem_1360;
  reg [31:0] _RAND_1360;
  reg [31:0] mem_1361;
  reg [31:0] _RAND_1361;
  reg [31:0] mem_1362;
  reg [31:0] _RAND_1362;
  reg [31:0] mem_1363;
  reg [31:0] _RAND_1363;
  reg [31:0] mem_1364;
  reg [31:0] _RAND_1364;
  reg [31:0] mem_1365;
  reg [31:0] _RAND_1365;
  reg [31:0] mem_1366;
  reg [31:0] _RAND_1366;
  reg [31:0] mem_1367;
  reg [31:0] _RAND_1367;
  reg [31:0] mem_1368;
  reg [31:0] _RAND_1368;
  reg [31:0] mem_1369;
  reg [31:0] _RAND_1369;
  reg [31:0] mem_1370;
  reg [31:0] _RAND_1370;
  reg [31:0] mem_1371;
  reg [31:0] _RAND_1371;
  reg [31:0] mem_1372;
  reg [31:0] _RAND_1372;
  reg [31:0] mem_1373;
  reg [31:0] _RAND_1373;
  reg [31:0] mem_1374;
  reg [31:0] _RAND_1374;
  reg [31:0] mem_1375;
  reg [31:0] _RAND_1375;
  reg [31:0] mem_1376;
  reg [31:0] _RAND_1376;
  reg [31:0] mem_1377;
  reg [31:0] _RAND_1377;
  reg [31:0] mem_1378;
  reg [31:0] _RAND_1378;
  reg [31:0] mem_1379;
  reg [31:0] _RAND_1379;
  reg [31:0] mem_1380;
  reg [31:0] _RAND_1380;
  reg [31:0] mem_1381;
  reg [31:0] _RAND_1381;
  reg [31:0] mem_1382;
  reg [31:0] _RAND_1382;
  reg [31:0] mem_1383;
  reg [31:0] _RAND_1383;
  reg [31:0] mem_1384;
  reg [31:0] _RAND_1384;
  reg [31:0] mem_1385;
  reg [31:0] _RAND_1385;
  reg [31:0] mem_1386;
  reg [31:0] _RAND_1386;
  reg [31:0] mem_1387;
  reg [31:0] _RAND_1387;
  reg [31:0] mem_1388;
  reg [31:0] _RAND_1388;
  reg [31:0] mem_1389;
  reg [31:0] _RAND_1389;
  reg [31:0] mem_1390;
  reg [31:0] _RAND_1390;
  reg [31:0] mem_1391;
  reg [31:0] _RAND_1391;
  reg [31:0] mem_1392;
  reg [31:0] _RAND_1392;
  reg [31:0] mem_1393;
  reg [31:0] _RAND_1393;
  reg [31:0] mem_1394;
  reg [31:0] _RAND_1394;
  reg [31:0] mem_1395;
  reg [31:0] _RAND_1395;
  reg [31:0] mem_1396;
  reg [31:0] _RAND_1396;
  reg [31:0] mem_1397;
  reg [31:0] _RAND_1397;
  reg [31:0] mem_1398;
  reg [31:0] _RAND_1398;
  reg [31:0] mem_1399;
  reg [31:0] _RAND_1399;
  reg [31:0] mem_1400;
  reg [31:0] _RAND_1400;
  reg [31:0] mem_1401;
  reg [31:0] _RAND_1401;
  reg [31:0] mem_1402;
  reg [31:0] _RAND_1402;
  reg [31:0] mem_1403;
  reg [31:0] _RAND_1403;
  reg [31:0] mem_1404;
  reg [31:0] _RAND_1404;
  reg [31:0] mem_1405;
  reg [31:0] _RAND_1405;
  reg [31:0] mem_1406;
  reg [31:0] _RAND_1406;
  reg [31:0] mem_1407;
  reg [31:0] _RAND_1407;
  reg [31:0] mem_1408;
  reg [31:0] _RAND_1408;
  reg [31:0] mem_1409;
  reg [31:0] _RAND_1409;
  reg [31:0] mem_1410;
  reg [31:0] _RAND_1410;
  reg [31:0] mem_1411;
  reg [31:0] _RAND_1411;
  reg [31:0] mem_1412;
  reg [31:0] _RAND_1412;
  reg [31:0] mem_1413;
  reg [31:0] _RAND_1413;
  reg [31:0] mem_1414;
  reg [31:0] _RAND_1414;
  reg [31:0] mem_1415;
  reg [31:0] _RAND_1415;
  reg [31:0] mem_1416;
  reg [31:0] _RAND_1416;
  reg [31:0] mem_1417;
  reg [31:0] _RAND_1417;
  reg [31:0] mem_1418;
  reg [31:0] _RAND_1418;
  reg [31:0] mem_1419;
  reg [31:0] _RAND_1419;
  reg [31:0] mem_1420;
  reg [31:0] _RAND_1420;
  reg [31:0] mem_1421;
  reg [31:0] _RAND_1421;
  reg [31:0] mem_1422;
  reg [31:0] _RAND_1422;
  reg [31:0] mem_1423;
  reg [31:0] _RAND_1423;
  reg [31:0] mem_1424;
  reg [31:0] _RAND_1424;
  reg [31:0] mem_1425;
  reg [31:0] _RAND_1425;
  reg [31:0] mem_1426;
  reg [31:0] _RAND_1426;
  reg [31:0] mem_1427;
  reg [31:0] _RAND_1427;
  reg [31:0] mem_1428;
  reg [31:0] _RAND_1428;
  reg [31:0] mem_1429;
  reg [31:0] _RAND_1429;
  reg [31:0] mem_1430;
  reg [31:0] _RAND_1430;
  reg [31:0] mem_1431;
  reg [31:0] _RAND_1431;
  reg [31:0] mem_1432;
  reg [31:0] _RAND_1432;
  reg [31:0] mem_1433;
  reg [31:0] _RAND_1433;
  reg [31:0] mem_1434;
  reg [31:0] _RAND_1434;
  reg [31:0] mem_1435;
  reg [31:0] _RAND_1435;
  reg [31:0] mem_1436;
  reg [31:0] _RAND_1436;
  reg [31:0] mem_1437;
  reg [31:0] _RAND_1437;
  reg [31:0] mem_1438;
  reg [31:0] _RAND_1438;
  reg [31:0] mem_1439;
  reg [31:0] _RAND_1439;
  reg [31:0] mem_1440;
  reg [31:0] _RAND_1440;
  reg [31:0] mem_1441;
  reg [31:0] _RAND_1441;
  reg [31:0] mem_1442;
  reg [31:0] _RAND_1442;
  reg [31:0] mem_1443;
  reg [31:0] _RAND_1443;
  reg [31:0] mem_1444;
  reg [31:0] _RAND_1444;
  reg [31:0] mem_1445;
  reg [31:0] _RAND_1445;
  reg [31:0] mem_1446;
  reg [31:0] _RAND_1446;
  reg [31:0] mem_1447;
  reg [31:0] _RAND_1447;
  reg [31:0] mem_1448;
  reg [31:0] _RAND_1448;
  reg [31:0] mem_1449;
  reg [31:0] _RAND_1449;
  reg [31:0] mem_1450;
  reg [31:0] _RAND_1450;
  reg [31:0] mem_1451;
  reg [31:0] _RAND_1451;
  reg [31:0] mem_1452;
  reg [31:0] _RAND_1452;
  reg [31:0] mem_1453;
  reg [31:0] _RAND_1453;
  reg [31:0] mem_1454;
  reg [31:0] _RAND_1454;
  reg [31:0] mem_1455;
  reg [31:0] _RAND_1455;
  reg [31:0] mem_1456;
  reg [31:0] _RAND_1456;
  reg [31:0] mem_1457;
  reg [31:0] _RAND_1457;
  reg [31:0] mem_1458;
  reg [31:0] _RAND_1458;
  reg [31:0] mem_1459;
  reg [31:0] _RAND_1459;
  reg [31:0] mem_1460;
  reg [31:0] _RAND_1460;
  reg [31:0] mem_1461;
  reg [31:0] _RAND_1461;
  reg [31:0] mem_1462;
  reg [31:0] _RAND_1462;
  reg [31:0] mem_1463;
  reg [31:0] _RAND_1463;
  reg [31:0] mem_1464;
  reg [31:0] _RAND_1464;
  reg [31:0] mem_1465;
  reg [31:0] _RAND_1465;
  reg [31:0] mem_1466;
  reg [31:0] _RAND_1466;
  reg [31:0] mem_1467;
  reg [31:0] _RAND_1467;
  reg [31:0] mem_1468;
  reg [31:0] _RAND_1468;
  reg [31:0] mem_1469;
  reg [31:0] _RAND_1469;
  reg [31:0] mem_1470;
  reg [31:0] _RAND_1470;
  reg [31:0] mem_1471;
  reg [31:0] _RAND_1471;
  reg [31:0] mem_1472;
  reg [31:0] _RAND_1472;
  reg [31:0] mem_1473;
  reg [31:0] _RAND_1473;
  reg [31:0] mem_1474;
  reg [31:0] _RAND_1474;
  reg [31:0] mem_1475;
  reg [31:0] _RAND_1475;
  reg [31:0] mem_1476;
  reg [31:0] _RAND_1476;
  reg [31:0] mem_1477;
  reg [31:0] _RAND_1477;
  reg [31:0] mem_1478;
  reg [31:0] _RAND_1478;
  reg [31:0] mem_1479;
  reg [31:0] _RAND_1479;
  reg [31:0] mem_1480;
  reg [31:0] _RAND_1480;
  reg [31:0] mem_1481;
  reg [31:0] _RAND_1481;
  reg [31:0] mem_1482;
  reg [31:0] _RAND_1482;
  reg [31:0] mem_1483;
  reg [31:0] _RAND_1483;
  reg [31:0] mem_1484;
  reg [31:0] _RAND_1484;
  reg [31:0] mem_1485;
  reg [31:0] _RAND_1485;
  reg [31:0] mem_1486;
  reg [31:0] _RAND_1486;
  reg [31:0] mem_1487;
  reg [31:0] _RAND_1487;
  reg [31:0] mem_1488;
  reg [31:0] _RAND_1488;
  reg [31:0] mem_1489;
  reg [31:0] _RAND_1489;
  reg [31:0] mem_1490;
  reg [31:0] _RAND_1490;
  reg [31:0] mem_1491;
  reg [31:0] _RAND_1491;
  reg [31:0] mem_1492;
  reg [31:0] _RAND_1492;
  reg [31:0] mem_1493;
  reg [31:0] _RAND_1493;
  reg [31:0] mem_1494;
  reg [31:0] _RAND_1494;
  reg [31:0] mem_1495;
  reg [31:0] _RAND_1495;
  reg [31:0] mem_1496;
  reg [31:0] _RAND_1496;
  reg [31:0] mem_1497;
  reg [31:0] _RAND_1497;
  reg [31:0] mem_1498;
  reg [31:0] _RAND_1498;
  reg [31:0] mem_1499;
  reg [31:0] _RAND_1499;
  reg [31:0] mem_1500;
  reg [31:0] _RAND_1500;
  reg [31:0] mem_1501;
  reg [31:0] _RAND_1501;
  reg [31:0] mem_1502;
  reg [31:0] _RAND_1502;
  reg [31:0] mem_1503;
  reg [31:0] _RAND_1503;
  reg [31:0] mem_1504;
  reg [31:0] _RAND_1504;
  reg [31:0] mem_1505;
  reg [31:0] _RAND_1505;
  reg [31:0] mem_1506;
  reg [31:0] _RAND_1506;
  reg [31:0] mem_1507;
  reg [31:0] _RAND_1507;
  reg [31:0] mem_1508;
  reg [31:0] _RAND_1508;
  reg [31:0] mem_1509;
  reg [31:0] _RAND_1509;
  reg [31:0] mem_1510;
  reg [31:0] _RAND_1510;
  reg [31:0] mem_1511;
  reg [31:0] _RAND_1511;
  reg [31:0] mem_1512;
  reg [31:0] _RAND_1512;
  reg [31:0] mem_1513;
  reg [31:0] _RAND_1513;
  reg [31:0] mem_1514;
  reg [31:0] _RAND_1514;
  reg [31:0] mem_1515;
  reg [31:0] _RAND_1515;
  reg [31:0] mem_1516;
  reg [31:0] _RAND_1516;
  reg [31:0] mem_1517;
  reg [31:0] _RAND_1517;
  reg [31:0] mem_1518;
  reg [31:0] _RAND_1518;
  reg [31:0] mem_1519;
  reg [31:0] _RAND_1519;
  reg [31:0] mem_1520;
  reg [31:0] _RAND_1520;
  reg [31:0] mem_1521;
  reg [31:0] _RAND_1521;
  reg [31:0] mem_1522;
  reg [31:0] _RAND_1522;
  reg [31:0] mem_1523;
  reg [31:0] _RAND_1523;
  reg [31:0] mem_1524;
  reg [31:0] _RAND_1524;
  reg [31:0] mem_1525;
  reg [31:0] _RAND_1525;
  reg [31:0] mem_1526;
  reg [31:0] _RAND_1526;
  reg [31:0] mem_1527;
  reg [31:0] _RAND_1527;
  reg [31:0] mem_1528;
  reg [31:0] _RAND_1528;
  reg [31:0] mem_1529;
  reg [31:0] _RAND_1529;
  reg [31:0] mem_1530;
  reg [31:0] _RAND_1530;
  reg [31:0] mem_1531;
  reg [31:0] _RAND_1531;
  reg [31:0] mem_1532;
  reg [31:0] _RAND_1532;
  reg [31:0] mem_1533;
  reg [31:0] _RAND_1533;
  reg [31:0] mem_1534;
  reg [31:0] _RAND_1534;
  reg [31:0] mem_1535;
  reg [31:0] _RAND_1535;
  reg [31:0] mem_1536;
  reg [31:0] _RAND_1536;
  reg [31:0] mem_1537;
  reg [31:0] _RAND_1537;
  reg [31:0] mem_1538;
  reg [31:0] _RAND_1538;
  reg [31:0] mem_1539;
  reg [31:0] _RAND_1539;
  reg [31:0] mem_1540;
  reg [31:0] _RAND_1540;
  reg [31:0] mem_1541;
  reg [31:0] _RAND_1541;
  reg [31:0] mem_1542;
  reg [31:0] _RAND_1542;
  reg [31:0] mem_1543;
  reg [31:0] _RAND_1543;
  reg [31:0] mem_1544;
  reg [31:0] _RAND_1544;
  reg [31:0] mem_1545;
  reg [31:0] _RAND_1545;
  reg [31:0] mem_1546;
  reg [31:0] _RAND_1546;
  reg [31:0] mem_1547;
  reg [31:0] _RAND_1547;
  reg [31:0] mem_1548;
  reg [31:0] _RAND_1548;
  reg [31:0] mem_1549;
  reg [31:0] _RAND_1549;
  reg [31:0] mem_1550;
  reg [31:0] _RAND_1550;
  reg [31:0] mem_1551;
  reg [31:0] _RAND_1551;
  reg [31:0] mem_1552;
  reg [31:0] _RAND_1552;
  reg [31:0] mem_1553;
  reg [31:0] _RAND_1553;
  reg [31:0] mem_1554;
  reg [31:0] _RAND_1554;
  reg [31:0] mem_1555;
  reg [31:0] _RAND_1555;
  reg [31:0] mem_1556;
  reg [31:0] _RAND_1556;
  reg [31:0] mem_1557;
  reg [31:0] _RAND_1557;
  reg [31:0] mem_1558;
  reg [31:0] _RAND_1558;
  reg [31:0] mem_1559;
  reg [31:0] _RAND_1559;
  reg [31:0] mem_1560;
  reg [31:0] _RAND_1560;
  reg [31:0] mem_1561;
  reg [31:0] _RAND_1561;
  reg [31:0] mem_1562;
  reg [31:0] _RAND_1562;
  reg [31:0] mem_1563;
  reg [31:0] _RAND_1563;
  reg [31:0] mem_1564;
  reg [31:0] _RAND_1564;
  reg [31:0] mem_1565;
  reg [31:0] _RAND_1565;
  reg [31:0] mem_1566;
  reg [31:0] _RAND_1566;
  reg [31:0] mem_1567;
  reg [31:0] _RAND_1567;
  reg [31:0] mem_1568;
  reg [31:0] _RAND_1568;
  reg [31:0] mem_1569;
  reg [31:0] _RAND_1569;
  reg [31:0] mem_1570;
  reg [31:0] _RAND_1570;
  reg [31:0] mem_1571;
  reg [31:0] _RAND_1571;
  reg [31:0] mem_1572;
  reg [31:0] _RAND_1572;
  reg [31:0] mem_1573;
  reg [31:0] _RAND_1573;
  reg [31:0] mem_1574;
  reg [31:0] _RAND_1574;
  reg [31:0] mem_1575;
  reg [31:0] _RAND_1575;
  reg [31:0] mem_1576;
  reg [31:0] _RAND_1576;
  reg [31:0] mem_1577;
  reg [31:0] _RAND_1577;
  reg [31:0] mem_1578;
  reg [31:0] _RAND_1578;
  reg [31:0] mem_1579;
  reg [31:0] _RAND_1579;
  reg [31:0] mem_1580;
  reg [31:0] _RAND_1580;
  reg [31:0] mem_1581;
  reg [31:0] _RAND_1581;
  reg [31:0] mem_1582;
  reg [31:0] _RAND_1582;
  reg [31:0] mem_1583;
  reg [31:0] _RAND_1583;
  reg [31:0] mem_1584;
  reg [31:0] _RAND_1584;
  reg [31:0] mem_1585;
  reg [31:0] _RAND_1585;
  reg [31:0] mem_1586;
  reg [31:0] _RAND_1586;
  reg [31:0] mem_1587;
  reg [31:0] _RAND_1587;
  reg [31:0] mem_1588;
  reg [31:0] _RAND_1588;
  reg [31:0] mem_1589;
  reg [31:0] _RAND_1589;
  reg [31:0] mem_1590;
  reg [31:0] _RAND_1590;
  reg [31:0] mem_1591;
  reg [31:0] _RAND_1591;
  reg [31:0] mem_1592;
  reg [31:0] _RAND_1592;
  reg [31:0] mem_1593;
  reg [31:0] _RAND_1593;
  reg [31:0] mem_1594;
  reg [31:0] _RAND_1594;
  reg [31:0] mem_1595;
  reg [31:0] _RAND_1595;
  reg [31:0] mem_1596;
  reg [31:0] _RAND_1596;
  reg [31:0] mem_1597;
  reg [31:0] _RAND_1597;
  reg [31:0] mem_1598;
  reg [31:0] _RAND_1598;
  reg [31:0] mem_1599;
  reg [31:0] _RAND_1599;
  reg [31:0] mem_1600;
  reg [31:0] _RAND_1600;
  reg [31:0] mem_1601;
  reg [31:0] _RAND_1601;
  reg [31:0] mem_1602;
  reg [31:0] _RAND_1602;
  reg [31:0] mem_1603;
  reg [31:0] _RAND_1603;
  reg [31:0] mem_1604;
  reg [31:0] _RAND_1604;
  reg [31:0] mem_1605;
  reg [31:0] _RAND_1605;
  reg [31:0] mem_1606;
  reg [31:0] _RAND_1606;
  reg [31:0] mem_1607;
  reg [31:0] _RAND_1607;
  reg [31:0] mem_1608;
  reg [31:0] _RAND_1608;
  reg [31:0] mem_1609;
  reg [31:0] _RAND_1609;
  reg [31:0] mem_1610;
  reg [31:0] _RAND_1610;
  reg [31:0] mem_1611;
  reg [31:0] _RAND_1611;
  reg [31:0] mem_1612;
  reg [31:0] _RAND_1612;
  reg [31:0] mem_1613;
  reg [31:0] _RAND_1613;
  reg [31:0] mem_1614;
  reg [31:0] _RAND_1614;
  reg [31:0] mem_1615;
  reg [31:0] _RAND_1615;
  reg [31:0] mem_1616;
  reg [31:0] _RAND_1616;
  reg [31:0] mem_1617;
  reg [31:0] _RAND_1617;
  reg [31:0] mem_1618;
  reg [31:0] _RAND_1618;
  reg [31:0] mem_1619;
  reg [31:0] _RAND_1619;
  reg [31:0] mem_1620;
  reg [31:0] _RAND_1620;
  reg [31:0] mem_1621;
  reg [31:0] _RAND_1621;
  reg [31:0] mem_1622;
  reg [31:0] _RAND_1622;
  reg [31:0] mem_1623;
  reg [31:0] _RAND_1623;
  reg [31:0] mem_1624;
  reg [31:0] _RAND_1624;
  reg [31:0] mem_1625;
  reg [31:0] _RAND_1625;
  reg [31:0] mem_1626;
  reg [31:0] _RAND_1626;
  reg [31:0] mem_1627;
  reg [31:0] _RAND_1627;
  reg [31:0] mem_1628;
  reg [31:0] _RAND_1628;
  reg [31:0] mem_1629;
  reg [31:0] _RAND_1629;
  reg [31:0] mem_1630;
  reg [31:0] _RAND_1630;
  reg [31:0] mem_1631;
  reg [31:0] _RAND_1631;
  reg [31:0] mem_1632;
  reg [31:0] _RAND_1632;
  reg [31:0] mem_1633;
  reg [31:0] _RAND_1633;
  reg [31:0] mem_1634;
  reg [31:0] _RAND_1634;
  reg [31:0] mem_1635;
  reg [31:0] _RAND_1635;
  reg [31:0] mem_1636;
  reg [31:0] _RAND_1636;
  reg [31:0] mem_1637;
  reg [31:0] _RAND_1637;
  reg [31:0] mem_1638;
  reg [31:0] _RAND_1638;
  reg [31:0] mem_1639;
  reg [31:0] _RAND_1639;
  reg [31:0] mem_1640;
  reg [31:0] _RAND_1640;
  reg [31:0] mem_1641;
  reg [31:0] _RAND_1641;
  reg [31:0] mem_1642;
  reg [31:0] _RAND_1642;
  reg [31:0] mem_1643;
  reg [31:0] _RAND_1643;
  reg [31:0] mem_1644;
  reg [31:0] _RAND_1644;
  reg [31:0] mem_1645;
  reg [31:0] _RAND_1645;
  reg [31:0] mem_1646;
  reg [31:0] _RAND_1646;
  reg [31:0] mem_1647;
  reg [31:0] _RAND_1647;
  reg [31:0] mem_1648;
  reg [31:0] _RAND_1648;
  reg [31:0] mem_1649;
  reg [31:0] _RAND_1649;
  reg [31:0] mem_1650;
  reg [31:0] _RAND_1650;
  reg [31:0] mem_1651;
  reg [31:0] _RAND_1651;
  reg [31:0] mem_1652;
  reg [31:0] _RAND_1652;
  reg [31:0] mem_1653;
  reg [31:0] _RAND_1653;
  reg [31:0] mem_1654;
  reg [31:0] _RAND_1654;
  reg [31:0] mem_1655;
  reg [31:0] _RAND_1655;
  reg [31:0] mem_1656;
  reg [31:0] _RAND_1656;
  reg [31:0] mem_1657;
  reg [31:0] _RAND_1657;
  reg [31:0] mem_1658;
  reg [31:0] _RAND_1658;
  reg [31:0] mem_1659;
  reg [31:0] _RAND_1659;
  reg [31:0] mem_1660;
  reg [31:0] _RAND_1660;
  reg [31:0] mem_1661;
  reg [31:0] _RAND_1661;
  reg [31:0] mem_1662;
  reg [31:0] _RAND_1662;
  reg [31:0] mem_1663;
  reg [31:0] _RAND_1663;
  reg [31:0] mem_1664;
  reg [31:0] _RAND_1664;
  reg [31:0] mem_1665;
  reg [31:0] _RAND_1665;
  reg [31:0] mem_1666;
  reg [31:0] _RAND_1666;
  reg [31:0] mem_1667;
  reg [31:0] _RAND_1667;
  reg [31:0] mem_1668;
  reg [31:0] _RAND_1668;
  reg [31:0] mem_1669;
  reg [31:0] _RAND_1669;
  reg [31:0] mem_1670;
  reg [31:0] _RAND_1670;
  reg [31:0] mem_1671;
  reg [31:0] _RAND_1671;
  reg [31:0] mem_1672;
  reg [31:0] _RAND_1672;
  reg [31:0] mem_1673;
  reg [31:0] _RAND_1673;
  reg [31:0] mem_1674;
  reg [31:0] _RAND_1674;
  reg [31:0] mem_1675;
  reg [31:0] _RAND_1675;
  reg [31:0] mem_1676;
  reg [31:0] _RAND_1676;
  reg [31:0] mem_1677;
  reg [31:0] _RAND_1677;
  reg [31:0] mem_1678;
  reg [31:0] _RAND_1678;
  reg [31:0] mem_1679;
  reg [31:0] _RAND_1679;
  reg [31:0] mem_1680;
  reg [31:0] _RAND_1680;
  reg [31:0] mem_1681;
  reg [31:0] _RAND_1681;
  reg [31:0] mem_1682;
  reg [31:0] _RAND_1682;
  reg [31:0] mem_1683;
  reg [31:0] _RAND_1683;
  reg [31:0] mem_1684;
  reg [31:0] _RAND_1684;
  reg [31:0] mem_1685;
  reg [31:0] _RAND_1685;
  reg [31:0] mem_1686;
  reg [31:0] _RAND_1686;
  reg [31:0] mem_1687;
  reg [31:0] _RAND_1687;
  reg [31:0] mem_1688;
  reg [31:0] _RAND_1688;
  reg [31:0] mem_1689;
  reg [31:0] _RAND_1689;
  reg [31:0] mem_1690;
  reg [31:0] _RAND_1690;
  reg [31:0] mem_1691;
  reg [31:0] _RAND_1691;
  reg [31:0] mem_1692;
  reg [31:0] _RAND_1692;
  reg [31:0] mem_1693;
  reg [31:0] _RAND_1693;
  reg [31:0] mem_1694;
  reg [31:0] _RAND_1694;
  reg [31:0] mem_1695;
  reg [31:0] _RAND_1695;
  reg [31:0] mem_1696;
  reg [31:0] _RAND_1696;
  reg [31:0] mem_1697;
  reg [31:0] _RAND_1697;
  reg [31:0] mem_1698;
  reg [31:0] _RAND_1698;
  reg [31:0] mem_1699;
  reg [31:0] _RAND_1699;
  reg [31:0] mem_1700;
  reg [31:0] _RAND_1700;
  reg [31:0] mem_1701;
  reg [31:0] _RAND_1701;
  reg [31:0] mem_1702;
  reg [31:0] _RAND_1702;
  reg [31:0] mem_1703;
  reg [31:0] _RAND_1703;
  reg [31:0] mem_1704;
  reg [31:0] _RAND_1704;
  reg [31:0] mem_1705;
  reg [31:0] _RAND_1705;
  reg [31:0] mem_1706;
  reg [31:0] _RAND_1706;
  reg [31:0] mem_1707;
  reg [31:0] _RAND_1707;
  reg [31:0] mem_1708;
  reg [31:0] _RAND_1708;
  reg [31:0] mem_1709;
  reg [31:0] _RAND_1709;
  reg [31:0] mem_1710;
  reg [31:0] _RAND_1710;
  reg [31:0] mem_1711;
  reg [31:0] _RAND_1711;
  reg [31:0] mem_1712;
  reg [31:0] _RAND_1712;
  reg [31:0] mem_1713;
  reg [31:0] _RAND_1713;
  reg [31:0] mem_1714;
  reg [31:0] _RAND_1714;
  reg [31:0] mem_1715;
  reg [31:0] _RAND_1715;
  reg [31:0] mem_1716;
  reg [31:0] _RAND_1716;
  reg [31:0] mem_1717;
  reg [31:0] _RAND_1717;
  reg [31:0] mem_1718;
  reg [31:0] _RAND_1718;
  reg [31:0] mem_1719;
  reg [31:0] _RAND_1719;
  reg [31:0] mem_1720;
  reg [31:0] _RAND_1720;
  reg [31:0] mem_1721;
  reg [31:0] _RAND_1721;
  reg [31:0] mem_1722;
  reg [31:0] _RAND_1722;
  reg [31:0] mem_1723;
  reg [31:0] _RAND_1723;
  reg [31:0] mem_1724;
  reg [31:0] _RAND_1724;
  reg [31:0] mem_1725;
  reg [31:0] _RAND_1725;
  reg [31:0] mem_1726;
  reg [31:0] _RAND_1726;
  reg [31:0] mem_1727;
  reg [31:0] _RAND_1727;
  reg [31:0] mem_1728;
  reg [31:0] _RAND_1728;
  reg [31:0] mem_1729;
  reg [31:0] _RAND_1729;
  reg [31:0] mem_1730;
  reg [31:0] _RAND_1730;
  reg [31:0] mem_1731;
  reg [31:0] _RAND_1731;
  reg [31:0] mem_1732;
  reg [31:0] _RAND_1732;
  reg [31:0] mem_1733;
  reg [31:0] _RAND_1733;
  reg [31:0] mem_1734;
  reg [31:0] _RAND_1734;
  reg [31:0] mem_1735;
  reg [31:0] _RAND_1735;
  reg [31:0] mem_1736;
  reg [31:0] _RAND_1736;
  reg [31:0] mem_1737;
  reg [31:0] _RAND_1737;
  reg [31:0] mem_1738;
  reg [31:0] _RAND_1738;
  reg [31:0] mem_1739;
  reg [31:0] _RAND_1739;
  reg [31:0] mem_1740;
  reg [31:0] _RAND_1740;
  reg [31:0] mem_1741;
  reg [31:0] _RAND_1741;
  reg [31:0] mem_1742;
  reg [31:0] _RAND_1742;
  reg [31:0] mem_1743;
  reg [31:0] _RAND_1743;
  reg [31:0] mem_1744;
  reg [31:0] _RAND_1744;
  reg [31:0] mem_1745;
  reg [31:0] _RAND_1745;
  reg [31:0] mem_1746;
  reg [31:0] _RAND_1746;
  reg [31:0] mem_1747;
  reg [31:0] _RAND_1747;
  reg [31:0] mem_1748;
  reg [31:0] _RAND_1748;
  reg [31:0] mem_1749;
  reg [31:0] _RAND_1749;
  reg [31:0] mem_1750;
  reg [31:0] _RAND_1750;
  reg [31:0] mem_1751;
  reg [31:0] _RAND_1751;
  reg [31:0] mem_1752;
  reg [31:0] _RAND_1752;
  reg [31:0] mem_1753;
  reg [31:0] _RAND_1753;
  reg [31:0] mem_1754;
  reg [31:0] _RAND_1754;
  reg [31:0] mem_1755;
  reg [31:0] _RAND_1755;
  reg [31:0] mem_1756;
  reg [31:0] _RAND_1756;
  reg [31:0] mem_1757;
  reg [31:0] _RAND_1757;
  reg [31:0] mem_1758;
  reg [31:0] _RAND_1758;
  reg [31:0] mem_1759;
  reg [31:0] _RAND_1759;
  reg [31:0] mem_1760;
  reg [31:0] _RAND_1760;
  reg [31:0] mem_1761;
  reg [31:0] _RAND_1761;
  reg [31:0] mem_1762;
  reg [31:0] _RAND_1762;
  reg [31:0] mem_1763;
  reg [31:0] _RAND_1763;
  reg [31:0] mem_1764;
  reg [31:0] _RAND_1764;
  reg [31:0] mem_1765;
  reg [31:0] _RAND_1765;
  reg [31:0] mem_1766;
  reg [31:0] _RAND_1766;
  reg [31:0] mem_1767;
  reg [31:0] _RAND_1767;
  reg [31:0] mem_1768;
  reg [31:0] _RAND_1768;
  reg [31:0] mem_1769;
  reg [31:0] _RAND_1769;
  reg [31:0] mem_1770;
  reg [31:0] _RAND_1770;
  reg [31:0] mem_1771;
  reg [31:0] _RAND_1771;
  reg [31:0] mem_1772;
  reg [31:0] _RAND_1772;
  reg [31:0] mem_1773;
  reg [31:0] _RAND_1773;
  reg [31:0] mem_1774;
  reg [31:0] _RAND_1774;
  reg [31:0] mem_1775;
  reg [31:0] _RAND_1775;
  reg [31:0] mem_1776;
  reg [31:0] _RAND_1776;
  reg [31:0] mem_1777;
  reg [31:0] _RAND_1777;
  reg [31:0] mem_1778;
  reg [31:0] _RAND_1778;
  reg [31:0] mem_1779;
  reg [31:0] _RAND_1779;
  reg [31:0] mem_1780;
  reg [31:0] _RAND_1780;
  reg [31:0] mem_1781;
  reg [31:0] _RAND_1781;
  reg [31:0] mem_1782;
  reg [31:0] _RAND_1782;
  reg [31:0] mem_1783;
  reg [31:0] _RAND_1783;
  reg [31:0] mem_1784;
  reg [31:0] _RAND_1784;
  reg [31:0] mem_1785;
  reg [31:0] _RAND_1785;
  reg [31:0] mem_1786;
  reg [31:0] _RAND_1786;
  reg [31:0] mem_1787;
  reg [31:0] _RAND_1787;
  reg [31:0] mem_1788;
  reg [31:0] _RAND_1788;
  reg [31:0] mem_1789;
  reg [31:0] _RAND_1789;
  reg [31:0] mem_1790;
  reg [31:0] _RAND_1790;
  reg [31:0] mem_1791;
  reg [31:0] _RAND_1791;
  reg [31:0] mem_1792;
  reg [31:0] _RAND_1792;
  reg [31:0] mem_1793;
  reg [31:0] _RAND_1793;
  reg [31:0] mem_1794;
  reg [31:0] _RAND_1794;
  reg [31:0] mem_1795;
  reg [31:0] _RAND_1795;
  reg [31:0] mem_1796;
  reg [31:0] _RAND_1796;
  reg [31:0] mem_1797;
  reg [31:0] _RAND_1797;
  reg [31:0] mem_1798;
  reg [31:0] _RAND_1798;
  reg [31:0] mem_1799;
  reg [31:0] _RAND_1799;
  reg [31:0] mem_1800;
  reg [31:0] _RAND_1800;
  reg [31:0] mem_1801;
  reg [31:0] _RAND_1801;
  reg [31:0] mem_1802;
  reg [31:0] _RAND_1802;
  reg [31:0] mem_1803;
  reg [31:0] _RAND_1803;
  reg [31:0] mem_1804;
  reg [31:0] _RAND_1804;
  reg [31:0] mem_1805;
  reg [31:0] _RAND_1805;
  reg [31:0] mem_1806;
  reg [31:0] _RAND_1806;
  reg [31:0] mem_1807;
  reg [31:0] _RAND_1807;
  reg [31:0] mem_1808;
  reg [31:0] _RAND_1808;
  reg [31:0] mem_1809;
  reg [31:0] _RAND_1809;
  reg [31:0] mem_1810;
  reg [31:0] _RAND_1810;
  reg [31:0] mem_1811;
  reg [31:0] _RAND_1811;
  reg [31:0] mem_1812;
  reg [31:0] _RAND_1812;
  reg [31:0] mem_1813;
  reg [31:0] _RAND_1813;
  reg [31:0] mem_1814;
  reg [31:0] _RAND_1814;
  reg [31:0] mem_1815;
  reg [31:0] _RAND_1815;
  reg [31:0] mem_1816;
  reg [31:0] _RAND_1816;
  reg [31:0] mem_1817;
  reg [31:0] _RAND_1817;
  reg [31:0] mem_1818;
  reg [31:0] _RAND_1818;
  reg [31:0] mem_1819;
  reg [31:0] _RAND_1819;
  reg [31:0] mem_1820;
  reg [31:0] _RAND_1820;
  reg [31:0] mem_1821;
  reg [31:0] _RAND_1821;
  reg [31:0] mem_1822;
  reg [31:0] _RAND_1822;
  reg [31:0] mem_1823;
  reg [31:0] _RAND_1823;
  reg [31:0] mem_1824;
  reg [31:0] _RAND_1824;
  reg [31:0] mem_1825;
  reg [31:0] _RAND_1825;
  reg [31:0] mem_1826;
  reg [31:0] _RAND_1826;
  reg [31:0] mem_1827;
  reg [31:0] _RAND_1827;
  reg [31:0] mem_1828;
  reg [31:0] _RAND_1828;
  reg [31:0] mem_1829;
  reg [31:0] _RAND_1829;
  reg [31:0] mem_1830;
  reg [31:0] _RAND_1830;
  reg [31:0] mem_1831;
  reg [31:0] _RAND_1831;
  reg [31:0] mem_1832;
  reg [31:0] _RAND_1832;
  reg [31:0] mem_1833;
  reg [31:0] _RAND_1833;
  reg [31:0] mem_1834;
  reg [31:0] _RAND_1834;
  reg [31:0] mem_1835;
  reg [31:0] _RAND_1835;
  reg [31:0] mem_1836;
  reg [31:0] _RAND_1836;
  reg [31:0] mem_1837;
  reg [31:0] _RAND_1837;
  reg [31:0] mem_1838;
  reg [31:0] _RAND_1838;
  reg [31:0] mem_1839;
  reg [31:0] _RAND_1839;
  reg [31:0] mem_1840;
  reg [31:0] _RAND_1840;
  reg [31:0] mem_1841;
  reg [31:0] _RAND_1841;
  reg [31:0] mem_1842;
  reg [31:0] _RAND_1842;
  reg [31:0] mem_1843;
  reg [31:0] _RAND_1843;
  reg [31:0] mem_1844;
  reg [31:0] _RAND_1844;
  reg [31:0] mem_1845;
  reg [31:0] _RAND_1845;
  reg [31:0] mem_1846;
  reg [31:0] _RAND_1846;
  reg [31:0] mem_1847;
  reg [31:0] _RAND_1847;
  reg [31:0] mem_1848;
  reg [31:0] _RAND_1848;
  reg [31:0] mem_1849;
  reg [31:0] _RAND_1849;
  reg [31:0] mem_1850;
  reg [31:0] _RAND_1850;
  reg [31:0] mem_1851;
  reg [31:0] _RAND_1851;
  reg [31:0] mem_1852;
  reg [31:0] _RAND_1852;
  reg [31:0] mem_1853;
  reg [31:0] _RAND_1853;
  reg [31:0] mem_1854;
  reg [31:0] _RAND_1854;
  reg [31:0] mem_1855;
  reg [31:0] _RAND_1855;
  reg [31:0] mem_1856;
  reg [31:0] _RAND_1856;
  reg [31:0] mem_1857;
  reg [31:0] _RAND_1857;
  reg [31:0] mem_1858;
  reg [31:0] _RAND_1858;
  reg [31:0] mem_1859;
  reg [31:0] _RAND_1859;
  reg [31:0] mem_1860;
  reg [31:0] _RAND_1860;
  reg [31:0] mem_1861;
  reg [31:0] _RAND_1861;
  reg [31:0] mem_1862;
  reg [31:0] _RAND_1862;
  reg [31:0] mem_1863;
  reg [31:0] _RAND_1863;
  reg [31:0] mem_1864;
  reg [31:0] _RAND_1864;
  reg [31:0] mem_1865;
  reg [31:0] _RAND_1865;
  reg [31:0] mem_1866;
  reg [31:0] _RAND_1866;
  reg [31:0] mem_1867;
  reg [31:0] _RAND_1867;
  reg [31:0] mem_1868;
  reg [31:0] _RAND_1868;
  reg [31:0] mem_1869;
  reg [31:0] _RAND_1869;
  reg [31:0] mem_1870;
  reg [31:0] _RAND_1870;
  reg [31:0] mem_1871;
  reg [31:0] _RAND_1871;
  reg [31:0] mem_1872;
  reg [31:0] _RAND_1872;
  reg [31:0] mem_1873;
  reg [31:0] _RAND_1873;
  reg [31:0] mem_1874;
  reg [31:0] _RAND_1874;
  reg [31:0] mem_1875;
  reg [31:0] _RAND_1875;
  reg [31:0] mem_1876;
  reg [31:0] _RAND_1876;
  reg [31:0] mem_1877;
  reg [31:0] _RAND_1877;
  reg [31:0] mem_1878;
  reg [31:0] _RAND_1878;
  reg [31:0] mem_1879;
  reg [31:0] _RAND_1879;
  reg [31:0] mem_1880;
  reg [31:0] _RAND_1880;
  reg [31:0] mem_1881;
  reg [31:0] _RAND_1881;
  reg [31:0] mem_1882;
  reg [31:0] _RAND_1882;
  reg [31:0] mem_1883;
  reg [31:0] _RAND_1883;
  reg [31:0] mem_1884;
  reg [31:0] _RAND_1884;
  reg [31:0] mem_1885;
  reg [31:0] _RAND_1885;
  reg [31:0] mem_1886;
  reg [31:0] _RAND_1886;
  reg [31:0] mem_1887;
  reg [31:0] _RAND_1887;
  reg [31:0] mem_1888;
  reg [31:0] _RAND_1888;
  reg [31:0] mem_1889;
  reg [31:0] _RAND_1889;
  reg [31:0] mem_1890;
  reg [31:0] _RAND_1890;
  reg [31:0] mem_1891;
  reg [31:0] _RAND_1891;
  reg [31:0] mem_1892;
  reg [31:0] _RAND_1892;
  reg [31:0] mem_1893;
  reg [31:0] _RAND_1893;
  reg [31:0] mem_1894;
  reg [31:0] _RAND_1894;
  reg [31:0] mem_1895;
  reg [31:0] _RAND_1895;
  reg [31:0] mem_1896;
  reg [31:0] _RAND_1896;
  reg [31:0] mem_1897;
  reg [31:0] _RAND_1897;
  reg [31:0] mem_1898;
  reg [31:0] _RAND_1898;
  reg [31:0] mem_1899;
  reg [31:0] _RAND_1899;
  reg [31:0] mem_1900;
  reg [31:0] _RAND_1900;
  reg [31:0] mem_1901;
  reg [31:0] _RAND_1901;
  reg [31:0] mem_1902;
  reg [31:0] _RAND_1902;
  reg [31:0] mem_1903;
  reg [31:0] _RAND_1903;
  reg [31:0] mem_1904;
  reg [31:0] _RAND_1904;
  reg [31:0] mem_1905;
  reg [31:0] _RAND_1905;
  reg [31:0] mem_1906;
  reg [31:0] _RAND_1906;
  reg [31:0] mem_1907;
  reg [31:0] _RAND_1907;
  reg [31:0] mem_1908;
  reg [31:0] _RAND_1908;
  reg [31:0] mem_1909;
  reg [31:0] _RAND_1909;
  reg [31:0] mem_1910;
  reg [31:0] _RAND_1910;
  reg [31:0] mem_1911;
  reg [31:0] _RAND_1911;
  reg [31:0] mem_1912;
  reg [31:0] _RAND_1912;
  reg [31:0] mem_1913;
  reg [31:0] _RAND_1913;
  reg [31:0] mem_1914;
  reg [31:0] _RAND_1914;
  reg [31:0] mem_1915;
  reg [31:0] _RAND_1915;
  reg [31:0] mem_1916;
  reg [31:0] _RAND_1916;
  reg [31:0] mem_1917;
  reg [31:0] _RAND_1917;
  reg [31:0] mem_1918;
  reg [31:0] _RAND_1918;
  reg [31:0] mem_1919;
  reg [31:0] _RAND_1919;
  reg [31:0] mem_1920;
  reg [31:0] _RAND_1920;
  reg [31:0] mem_1921;
  reg [31:0] _RAND_1921;
  reg [31:0] mem_1922;
  reg [31:0] _RAND_1922;
  reg [31:0] mem_1923;
  reg [31:0] _RAND_1923;
  reg [31:0] mem_1924;
  reg [31:0] _RAND_1924;
  reg [31:0] mem_1925;
  reg [31:0] _RAND_1925;
  reg [31:0] mem_1926;
  reg [31:0] _RAND_1926;
  reg [31:0] mem_1927;
  reg [31:0] _RAND_1927;
  reg [31:0] mem_1928;
  reg [31:0] _RAND_1928;
  reg [31:0] mem_1929;
  reg [31:0] _RAND_1929;
  reg [31:0] mem_1930;
  reg [31:0] _RAND_1930;
  reg [31:0] mem_1931;
  reg [31:0] _RAND_1931;
  reg [31:0] mem_1932;
  reg [31:0] _RAND_1932;
  reg [31:0] mem_1933;
  reg [31:0] _RAND_1933;
  reg [31:0] mem_1934;
  reg [31:0] _RAND_1934;
  reg [31:0] mem_1935;
  reg [31:0] _RAND_1935;
  reg [31:0] mem_1936;
  reg [31:0] _RAND_1936;
  reg [31:0] mem_1937;
  reg [31:0] _RAND_1937;
  reg [31:0] mem_1938;
  reg [31:0] _RAND_1938;
  reg [31:0] mem_1939;
  reg [31:0] _RAND_1939;
  reg [31:0] mem_1940;
  reg [31:0] _RAND_1940;
  reg [31:0] mem_1941;
  reg [31:0] _RAND_1941;
  reg [31:0] mem_1942;
  reg [31:0] _RAND_1942;
  reg [31:0] mem_1943;
  reg [31:0] _RAND_1943;
  reg [31:0] mem_1944;
  reg [31:0] _RAND_1944;
  reg [31:0] mem_1945;
  reg [31:0] _RAND_1945;
  reg [31:0] mem_1946;
  reg [31:0] _RAND_1946;
  reg [31:0] mem_1947;
  reg [31:0] _RAND_1947;
  reg [31:0] mem_1948;
  reg [31:0] _RAND_1948;
  reg [31:0] mem_1949;
  reg [31:0] _RAND_1949;
  reg [31:0] mem_1950;
  reg [31:0] _RAND_1950;
  reg [31:0] mem_1951;
  reg [31:0] _RAND_1951;
  reg [31:0] mem_1952;
  reg [31:0] _RAND_1952;
  reg [31:0] mem_1953;
  reg [31:0] _RAND_1953;
  reg [31:0] mem_1954;
  reg [31:0] _RAND_1954;
  reg [31:0] mem_1955;
  reg [31:0] _RAND_1955;
  reg [31:0] mem_1956;
  reg [31:0] _RAND_1956;
  reg [31:0] mem_1957;
  reg [31:0] _RAND_1957;
  reg [31:0] mem_1958;
  reg [31:0] _RAND_1958;
  reg [31:0] mem_1959;
  reg [31:0] _RAND_1959;
  reg [31:0] mem_1960;
  reg [31:0] _RAND_1960;
  reg [31:0] mem_1961;
  reg [31:0] _RAND_1961;
  reg [31:0] mem_1962;
  reg [31:0] _RAND_1962;
  reg [31:0] mem_1963;
  reg [31:0] _RAND_1963;
  reg [31:0] mem_1964;
  reg [31:0] _RAND_1964;
  reg [31:0] mem_1965;
  reg [31:0] _RAND_1965;
  reg [31:0] mem_1966;
  reg [31:0] _RAND_1966;
  reg [31:0] mem_1967;
  reg [31:0] _RAND_1967;
  reg [31:0] mem_1968;
  reg [31:0] _RAND_1968;
  reg [31:0] mem_1969;
  reg [31:0] _RAND_1969;
  reg [31:0] mem_1970;
  reg [31:0] _RAND_1970;
  reg [31:0] mem_1971;
  reg [31:0] _RAND_1971;
  reg [31:0] mem_1972;
  reg [31:0] _RAND_1972;
  reg [31:0] mem_1973;
  reg [31:0] _RAND_1973;
  reg [31:0] mem_1974;
  reg [31:0] _RAND_1974;
  reg [31:0] mem_1975;
  reg [31:0] _RAND_1975;
  reg [31:0] mem_1976;
  reg [31:0] _RAND_1976;
  reg [31:0] mem_1977;
  reg [31:0] _RAND_1977;
  reg [31:0] mem_1978;
  reg [31:0] _RAND_1978;
  reg [31:0] mem_1979;
  reg [31:0] _RAND_1979;
  reg [31:0] mem_1980;
  reg [31:0] _RAND_1980;
  reg [31:0] mem_1981;
  reg [31:0] _RAND_1981;
  reg [31:0] mem_1982;
  reg [31:0] _RAND_1982;
  reg [31:0] mem_1983;
  reg [31:0] _RAND_1983;
  reg [31:0] mem_1984;
  reg [31:0] _RAND_1984;
  reg [31:0] mem_1985;
  reg [31:0] _RAND_1985;
  reg [31:0] mem_1986;
  reg [31:0] _RAND_1986;
  reg [31:0] mem_1987;
  reg [31:0] _RAND_1987;
  reg [31:0] mem_1988;
  reg [31:0] _RAND_1988;
  reg [31:0] mem_1989;
  reg [31:0] _RAND_1989;
  reg [31:0] mem_1990;
  reg [31:0] _RAND_1990;
  reg [31:0] mem_1991;
  reg [31:0] _RAND_1991;
  reg [31:0] mem_1992;
  reg [31:0] _RAND_1992;
  reg [31:0] mem_1993;
  reg [31:0] _RAND_1993;
  reg [31:0] mem_1994;
  reg [31:0] _RAND_1994;
  reg [31:0] mem_1995;
  reg [31:0] _RAND_1995;
  reg [31:0] mem_1996;
  reg [31:0] _RAND_1996;
  reg [31:0] mem_1997;
  reg [31:0] _RAND_1997;
  reg [31:0] mem_1998;
  reg [31:0] _RAND_1998;
  reg [31:0] mem_1999;
  reg [31:0] _RAND_1999;
  reg [31:0] mem_2000;
  reg [31:0] _RAND_2000;
  reg [31:0] mem_2001;
  reg [31:0] _RAND_2001;
  reg [31:0] mem_2002;
  reg [31:0] _RAND_2002;
  reg [31:0] mem_2003;
  reg [31:0] _RAND_2003;
  reg [31:0] mem_2004;
  reg [31:0] _RAND_2004;
  reg [31:0] mem_2005;
  reg [31:0] _RAND_2005;
  reg [31:0] mem_2006;
  reg [31:0] _RAND_2006;
  reg [31:0] mem_2007;
  reg [31:0] _RAND_2007;
  reg [31:0] mem_2008;
  reg [31:0] _RAND_2008;
  reg [31:0] mem_2009;
  reg [31:0] _RAND_2009;
  reg [31:0] mem_2010;
  reg [31:0] _RAND_2010;
  reg [31:0] mem_2011;
  reg [31:0] _RAND_2011;
  reg [31:0] mem_2012;
  reg [31:0] _RAND_2012;
  reg [31:0] mem_2013;
  reg [31:0] _RAND_2013;
  reg [31:0] mem_2014;
  reg [31:0] _RAND_2014;
  reg [31:0] mem_2015;
  reg [31:0] _RAND_2015;
  reg [31:0] mem_2016;
  reg [31:0] _RAND_2016;
  reg [31:0] mem_2017;
  reg [31:0] _RAND_2017;
  reg [31:0] mem_2018;
  reg [31:0] _RAND_2018;
  reg [31:0] mem_2019;
  reg [31:0] _RAND_2019;
  reg [31:0] mem_2020;
  reg [31:0] _RAND_2020;
  reg [31:0] mem_2021;
  reg [31:0] _RAND_2021;
  reg [31:0] mem_2022;
  reg [31:0] _RAND_2022;
  reg [31:0] mem_2023;
  reg [31:0] _RAND_2023;
  reg [31:0] mem_2024;
  reg [31:0] _RAND_2024;
  reg [31:0] mem_2025;
  reg [31:0] _RAND_2025;
  reg [31:0] mem_2026;
  reg [31:0] _RAND_2026;
  reg [31:0] mem_2027;
  reg [31:0] _RAND_2027;
  reg [31:0] mem_2028;
  reg [31:0] _RAND_2028;
  reg [31:0] mem_2029;
  reg [31:0] _RAND_2029;
  reg [31:0] mem_2030;
  reg [31:0] _RAND_2030;
  reg [31:0] mem_2031;
  reg [31:0] _RAND_2031;
  reg [31:0] mem_2032;
  reg [31:0] _RAND_2032;
  reg [31:0] mem_2033;
  reg [31:0] _RAND_2033;
  reg [31:0] mem_2034;
  reg [31:0] _RAND_2034;
  reg [31:0] mem_2035;
  reg [31:0] _RAND_2035;
  reg [31:0] mem_2036;
  reg [31:0] _RAND_2036;
  reg [31:0] mem_2037;
  reg [31:0] _RAND_2037;
  reg [31:0] mem_2038;
  reg [31:0] _RAND_2038;
  reg [31:0] mem_2039;
  reg [31:0] _RAND_2039;
  reg [31:0] mem_2040;
  reg [31:0] _RAND_2040;
  reg [31:0] mem_2041;
  reg [31:0] _RAND_2041;
  reg [31:0] mem_2042;
  reg [31:0] _RAND_2042;
  reg [31:0] mem_2043;
  reg [31:0] _RAND_2043;
  reg [31:0] mem_2044;
  reg [31:0] _RAND_2044;
  reg [31:0] mem_2045;
  reg [31:0] _RAND_2045;
  reg [31:0] mem_2046;
  reg [31:0] _RAND_2046;
  reg [31:0] mem_2047;
  reg [31:0] _RAND_2047;
  wire [7:0] toWrite_0;
  wire [7:0] toWrite_1;
  wire [7:0] toWrite_2;
  wire [7:0] toWrite_3;
  wire  _T_12316;
  wire [7:0] _T_12319;
  wire [10:0] _T_12323;
  wire [31:0] _GEN_0;
  wire [31:0] _GEN_6;
  wire [31:0] _GEN_7;
  wire [31:0] _GEN_8;
  wire [31:0] _GEN_9;
  wire [31:0] _GEN_10;
  wire [31:0] _GEN_11;
  wire [31:0] _GEN_12;
  wire [31:0] _GEN_13;
  wire [31:0] _GEN_14;
  wire [31:0] _GEN_15;
  wire [31:0] _GEN_16;
  wire [31:0] _GEN_17;
  wire [31:0] _GEN_18;
  wire [31:0] _GEN_19;
  wire [31:0] _GEN_20;
  wire [31:0] _GEN_21;
  wire [31:0] _GEN_22;
  wire [31:0] _GEN_23;
  wire [31:0] _GEN_24;
  wire [31:0] _GEN_25;
  wire [31:0] _GEN_26;
  wire [31:0] _GEN_27;
  wire [31:0] _GEN_28;
  wire [31:0] _GEN_29;
  wire [31:0] _GEN_30;
  wire [31:0] _GEN_31;
  wire [31:0] _GEN_32;
  wire [31:0] _GEN_33;
  wire [31:0] _GEN_34;
  wire [31:0] _GEN_35;
  wire [31:0] _GEN_36;
  wire [31:0] _GEN_37;
  wire [31:0] _GEN_38;
  wire [31:0] _GEN_39;
  wire [31:0] _GEN_40;
  wire [31:0] _GEN_41;
  wire [31:0] _GEN_42;
  wire [31:0] _GEN_43;
  wire [31:0] _GEN_44;
  wire [31:0] _GEN_45;
  wire [31:0] _GEN_46;
  wire [31:0] _GEN_47;
  wire [31:0] _GEN_48;
  wire [31:0] _GEN_49;
  wire [31:0] _GEN_50;
  wire [31:0] _GEN_51;
  wire [31:0] _GEN_52;
  wire [31:0] _GEN_53;
  wire [31:0] _GEN_54;
  wire [31:0] _GEN_55;
  wire [31:0] _GEN_56;
  wire [31:0] _GEN_57;
  wire [31:0] _GEN_58;
  wire [31:0] _GEN_59;
  wire [31:0] _GEN_60;
  wire [31:0] _GEN_61;
  wire [31:0] _GEN_62;
  wire [31:0] _GEN_63;
  wire [31:0] _GEN_64;
  wire [31:0] _GEN_65;
  wire [31:0] _GEN_66;
  wire [31:0] _GEN_67;
  wire [31:0] _GEN_68;
  wire [31:0] _GEN_69;
  wire [31:0] _GEN_70;
  wire [31:0] _GEN_71;
  wire [31:0] _GEN_72;
  wire [31:0] _GEN_73;
  wire [31:0] _GEN_74;
  wire [31:0] _GEN_75;
  wire [31:0] _GEN_76;
  wire [31:0] _GEN_77;
  wire [31:0] _GEN_78;
  wire [31:0] _GEN_79;
  wire [31:0] _GEN_80;
  wire [31:0] _GEN_81;
  wire [31:0] _GEN_82;
  wire [31:0] _GEN_83;
  wire [31:0] _GEN_84;
  wire [31:0] _GEN_85;
  wire [31:0] _GEN_86;
  wire [31:0] _GEN_87;
  wire [31:0] _GEN_88;
  wire [31:0] _GEN_89;
  wire [31:0] _GEN_90;
  wire [31:0] _GEN_91;
  wire [31:0] _GEN_92;
  wire [31:0] _GEN_93;
  wire [31:0] _GEN_94;
  wire [31:0] _GEN_95;
  wire [31:0] _GEN_96;
  wire [31:0] _GEN_97;
  wire [31:0] _GEN_98;
  wire [31:0] _GEN_99;
  wire [31:0] _GEN_100;
  wire [31:0] _GEN_101;
  wire [31:0] _GEN_102;
  wire [31:0] _GEN_103;
  wire [31:0] _GEN_104;
  wire [31:0] _GEN_105;
  wire [31:0] _GEN_106;
  wire [31:0] _GEN_107;
  wire [31:0] _GEN_108;
  wire [31:0] _GEN_109;
  wire [31:0] _GEN_110;
  wire [31:0] _GEN_111;
  wire [31:0] _GEN_112;
  wire [31:0] _GEN_113;
  wire [31:0] _GEN_114;
  wire [31:0] _GEN_115;
  wire [31:0] _GEN_116;
  wire [31:0] _GEN_117;
  wire [31:0] _GEN_118;
  wire [31:0] _GEN_119;
  wire [31:0] _GEN_120;
  wire [31:0] _GEN_121;
  wire [31:0] _GEN_122;
  wire [31:0] _GEN_123;
  wire [31:0] _GEN_124;
  wire [31:0] _GEN_125;
  wire [31:0] _GEN_126;
  wire [31:0] _GEN_127;
  wire [31:0] _GEN_128;
  wire [31:0] _GEN_129;
  wire [31:0] _GEN_130;
  wire [31:0] _GEN_131;
  wire [31:0] _GEN_132;
  wire [31:0] _GEN_133;
  wire [31:0] _GEN_134;
  wire [31:0] _GEN_135;
  wire [31:0] _GEN_136;
  wire [31:0] _GEN_137;
  wire [31:0] _GEN_138;
  wire [31:0] _GEN_139;
  wire [31:0] _GEN_140;
  wire [31:0] _GEN_141;
  wire [31:0] _GEN_142;
  wire [31:0] _GEN_143;
  wire [31:0] _GEN_144;
  wire [31:0] _GEN_145;
  wire [31:0] _GEN_146;
  wire [31:0] _GEN_147;
  wire [31:0] _GEN_148;
  wire [31:0] _GEN_149;
  wire [31:0] _GEN_150;
  wire [31:0] _GEN_151;
  wire [31:0] _GEN_152;
  wire [31:0] _GEN_153;
  wire [31:0] _GEN_154;
  wire [31:0] _GEN_155;
  wire [31:0] _GEN_156;
  wire [31:0] _GEN_157;
  wire [31:0] _GEN_158;
  wire [31:0] _GEN_159;
  wire [31:0] _GEN_160;
  wire [31:0] _GEN_161;
  wire [31:0] _GEN_162;
  wire [31:0] _GEN_163;
  wire [31:0] _GEN_164;
  wire [31:0] _GEN_165;
  wire [31:0] _GEN_166;
  wire [31:0] _GEN_167;
  wire [31:0] _GEN_168;
  wire [31:0] _GEN_169;
  wire [31:0] _GEN_170;
  wire [31:0] _GEN_171;
  wire [31:0] _GEN_172;
  wire [31:0] _GEN_173;
  wire [31:0] _GEN_174;
  wire [31:0] _GEN_175;
  wire [31:0] _GEN_176;
  wire [31:0] _GEN_177;
  wire [31:0] _GEN_178;
  wire [31:0] _GEN_179;
  wire [31:0] _GEN_180;
  wire [31:0] _GEN_181;
  wire [31:0] _GEN_182;
  wire [31:0] _GEN_183;
  wire [31:0] _GEN_184;
  wire [31:0] _GEN_185;
  wire [31:0] _GEN_186;
  wire [31:0] _GEN_187;
  wire [31:0] _GEN_188;
  wire [31:0] _GEN_189;
  wire [31:0] _GEN_190;
  wire [31:0] _GEN_191;
  wire [31:0] _GEN_192;
  wire [31:0] _GEN_193;
  wire [31:0] _GEN_194;
  wire [31:0] _GEN_195;
  wire [31:0] _GEN_196;
  wire [31:0] _GEN_197;
  wire [31:0] _GEN_198;
  wire [31:0] _GEN_199;
  wire [31:0] _GEN_200;
  wire [31:0] _GEN_201;
  wire [31:0] _GEN_202;
  wire [31:0] _GEN_203;
  wire [31:0] _GEN_204;
  wire [31:0] _GEN_205;
  wire [31:0] _GEN_206;
  wire [31:0] _GEN_207;
  wire [31:0] _GEN_208;
  wire [31:0] _GEN_209;
  wire [31:0] _GEN_210;
  wire [31:0] _GEN_211;
  wire [31:0] _GEN_212;
  wire [31:0] _GEN_213;
  wire [31:0] _GEN_214;
  wire [31:0] _GEN_215;
  wire [31:0] _GEN_216;
  wire [31:0] _GEN_217;
  wire [31:0] _GEN_218;
  wire [31:0] _GEN_219;
  wire [31:0] _GEN_220;
  wire [31:0] _GEN_221;
  wire [31:0] _GEN_222;
  wire [31:0] _GEN_223;
  wire [31:0] _GEN_224;
  wire [31:0] _GEN_225;
  wire [31:0] _GEN_226;
  wire [31:0] _GEN_227;
  wire [31:0] _GEN_228;
  wire [31:0] _GEN_229;
  wire [31:0] _GEN_230;
  wire [31:0] _GEN_231;
  wire [31:0] _GEN_232;
  wire [31:0] _GEN_233;
  wire [31:0] _GEN_234;
  wire [31:0] _GEN_235;
  wire [31:0] _GEN_236;
  wire [31:0] _GEN_237;
  wire [31:0] _GEN_238;
  wire [31:0] _GEN_239;
  wire [31:0] _GEN_240;
  wire [31:0] _GEN_241;
  wire [31:0] _GEN_242;
  wire [31:0] _GEN_243;
  wire [31:0] _GEN_244;
  wire [31:0] _GEN_245;
  wire [31:0] _GEN_246;
  wire [31:0] _GEN_247;
  wire [31:0] _GEN_248;
  wire [31:0] _GEN_249;
  wire [31:0] _GEN_250;
  wire [31:0] _GEN_251;
  wire [31:0] _GEN_252;
  wire [31:0] _GEN_253;
  wire [31:0] _GEN_254;
  wire [31:0] _GEN_255;
  wire [31:0] _GEN_256;
  wire [31:0] _GEN_257;
  wire [31:0] _GEN_258;
  wire [31:0] _GEN_259;
  wire [31:0] _GEN_260;
  wire [31:0] _GEN_261;
  wire [31:0] _GEN_262;
  wire [31:0] _GEN_263;
  wire [31:0] _GEN_264;
  wire [31:0] _GEN_265;
  wire [31:0] _GEN_266;
  wire [31:0] _GEN_267;
  wire [31:0] _GEN_268;
  wire [31:0] _GEN_269;
  wire [31:0] _GEN_270;
  wire [31:0] _GEN_271;
  wire [31:0] _GEN_272;
  wire [31:0] _GEN_273;
  wire [31:0] _GEN_274;
  wire [31:0] _GEN_275;
  wire [31:0] _GEN_276;
  wire [31:0] _GEN_277;
  wire [31:0] _GEN_278;
  wire [31:0] _GEN_279;
  wire [31:0] _GEN_280;
  wire [31:0] _GEN_281;
  wire [31:0] _GEN_282;
  wire [31:0] _GEN_283;
  wire [31:0] _GEN_284;
  wire [31:0] _GEN_285;
  wire [31:0] _GEN_286;
  wire [31:0] _GEN_287;
  wire [31:0] _GEN_288;
  wire [31:0] _GEN_289;
  wire [31:0] _GEN_290;
  wire [31:0] _GEN_291;
  wire [31:0] _GEN_292;
  wire [31:0] _GEN_293;
  wire [31:0] _GEN_294;
  wire [31:0] _GEN_295;
  wire [31:0] _GEN_296;
  wire [31:0] _GEN_297;
  wire [31:0] _GEN_298;
  wire [31:0] _GEN_299;
  wire [31:0] _GEN_300;
  wire [31:0] _GEN_301;
  wire [31:0] _GEN_302;
  wire [31:0] _GEN_303;
  wire [31:0] _GEN_304;
  wire [31:0] _GEN_305;
  wire [31:0] _GEN_306;
  wire [31:0] _GEN_307;
  wire [31:0] _GEN_308;
  wire [31:0] _GEN_309;
  wire [31:0] _GEN_310;
  wire [31:0] _GEN_311;
  wire [31:0] _GEN_312;
  wire [31:0] _GEN_313;
  wire [31:0] _GEN_314;
  wire [31:0] _GEN_315;
  wire [31:0] _GEN_316;
  wire [31:0] _GEN_317;
  wire [31:0] _GEN_318;
  wire [31:0] _GEN_319;
  wire [31:0] _GEN_320;
  wire [31:0] _GEN_321;
  wire [31:0] _GEN_322;
  wire [31:0] _GEN_323;
  wire [31:0] _GEN_324;
  wire [31:0] _GEN_325;
  wire [31:0] _GEN_326;
  wire [31:0] _GEN_327;
  wire [31:0] _GEN_328;
  wire [31:0] _GEN_329;
  wire [31:0] _GEN_330;
  wire [31:0] _GEN_331;
  wire [31:0] _GEN_332;
  wire [31:0] _GEN_333;
  wire [31:0] _GEN_334;
  wire [31:0] _GEN_335;
  wire [31:0] _GEN_336;
  wire [31:0] _GEN_337;
  wire [31:0] _GEN_338;
  wire [31:0] _GEN_339;
  wire [31:0] _GEN_340;
  wire [31:0] _GEN_341;
  wire [31:0] _GEN_342;
  wire [31:0] _GEN_343;
  wire [31:0] _GEN_344;
  wire [31:0] _GEN_345;
  wire [31:0] _GEN_346;
  wire [31:0] _GEN_347;
  wire [31:0] _GEN_348;
  wire [31:0] _GEN_349;
  wire [31:0] _GEN_350;
  wire [31:0] _GEN_351;
  wire [31:0] _GEN_352;
  wire [31:0] _GEN_353;
  wire [31:0] _GEN_354;
  wire [31:0] _GEN_355;
  wire [31:0] _GEN_356;
  wire [31:0] _GEN_357;
  wire [31:0] _GEN_358;
  wire [31:0] _GEN_359;
  wire [31:0] _GEN_360;
  wire [31:0] _GEN_361;
  wire [31:0] _GEN_362;
  wire [31:0] _GEN_363;
  wire [31:0] _GEN_364;
  wire [31:0] _GEN_365;
  wire [31:0] _GEN_366;
  wire [31:0] _GEN_367;
  wire [31:0] _GEN_368;
  wire [31:0] _GEN_369;
  wire [31:0] _GEN_370;
  wire [31:0] _GEN_371;
  wire [31:0] _GEN_372;
  wire [31:0] _GEN_373;
  wire [31:0] _GEN_374;
  wire [31:0] _GEN_375;
  wire [31:0] _GEN_376;
  wire [31:0] _GEN_377;
  wire [31:0] _GEN_378;
  wire [31:0] _GEN_379;
  wire [31:0] _GEN_380;
  wire [31:0] _GEN_381;
  wire [31:0] _GEN_382;
  wire [31:0] _GEN_383;
  wire [31:0] _GEN_384;
  wire [31:0] _GEN_385;
  wire [31:0] _GEN_386;
  wire [31:0] _GEN_387;
  wire [31:0] _GEN_388;
  wire [31:0] _GEN_389;
  wire [31:0] _GEN_390;
  wire [31:0] _GEN_391;
  wire [31:0] _GEN_392;
  wire [31:0] _GEN_393;
  wire [31:0] _GEN_394;
  wire [31:0] _GEN_395;
  wire [31:0] _GEN_396;
  wire [31:0] _GEN_397;
  wire [31:0] _GEN_398;
  wire [31:0] _GEN_399;
  wire [31:0] _GEN_400;
  wire [31:0] _GEN_401;
  wire [31:0] _GEN_402;
  wire [31:0] _GEN_403;
  wire [31:0] _GEN_404;
  wire [31:0] _GEN_405;
  wire [31:0] _GEN_406;
  wire [31:0] _GEN_407;
  wire [31:0] _GEN_408;
  wire [31:0] _GEN_409;
  wire [31:0] _GEN_410;
  wire [31:0] _GEN_411;
  wire [31:0] _GEN_412;
  wire [31:0] _GEN_413;
  wire [31:0] _GEN_414;
  wire [31:0] _GEN_415;
  wire [31:0] _GEN_416;
  wire [31:0] _GEN_417;
  wire [31:0] _GEN_418;
  wire [31:0] _GEN_419;
  wire [31:0] _GEN_420;
  wire [31:0] _GEN_421;
  wire [31:0] _GEN_422;
  wire [31:0] _GEN_423;
  wire [31:0] _GEN_424;
  wire [31:0] _GEN_425;
  wire [31:0] _GEN_426;
  wire [31:0] _GEN_427;
  wire [31:0] _GEN_428;
  wire [31:0] _GEN_429;
  wire [31:0] _GEN_430;
  wire [31:0] _GEN_431;
  wire [31:0] _GEN_432;
  wire [31:0] _GEN_433;
  wire [31:0] _GEN_434;
  wire [31:0] _GEN_435;
  wire [31:0] _GEN_436;
  wire [31:0] _GEN_437;
  wire [31:0] _GEN_438;
  wire [31:0] _GEN_439;
  wire [31:0] _GEN_440;
  wire [31:0] _GEN_441;
  wire [31:0] _GEN_442;
  wire [31:0] _GEN_443;
  wire [31:0] _GEN_444;
  wire [31:0] _GEN_445;
  wire [31:0] _GEN_446;
  wire [31:0] _GEN_447;
  wire [31:0] _GEN_448;
  wire [31:0] _GEN_449;
  wire [31:0] _GEN_450;
  wire [31:0] _GEN_451;
  wire [31:0] _GEN_452;
  wire [31:0] _GEN_453;
  wire [31:0] _GEN_454;
  wire [31:0] _GEN_455;
  wire [31:0] _GEN_456;
  wire [31:0] _GEN_457;
  wire [31:0] _GEN_458;
  wire [31:0] _GEN_459;
  wire [31:0] _GEN_460;
  wire [31:0] _GEN_461;
  wire [31:0] _GEN_462;
  wire [31:0] _GEN_463;
  wire [31:0] _GEN_464;
  wire [31:0] _GEN_465;
  wire [31:0] _GEN_466;
  wire [31:0] _GEN_467;
  wire [31:0] _GEN_468;
  wire [31:0] _GEN_469;
  wire [31:0] _GEN_470;
  wire [31:0] _GEN_471;
  wire [31:0] _GEN_472;
  wire [31:0] _GEN_473;
  wire [31:0] _GEN_474;
  wire [31:0] _GEN_475;
  wire [31:0] _GEN_476;
  wire [31:0] _GEN_477;
  wire [31:0] _GEN_478;
  wire [31:0] _GEN_479;
  wire [31:0] _GEN_480;
  wire [31:0] _GEN_481;
  wire [31:0] _GEN_482;
  wire [31:0] _GEN_483;
  wire [31:0] _GEN_484;
  wire [31:0] _GEN_485;
  wire [31:0] _GEN_486;
  wire [31:0] _GEN_487;
  wire [31:0] _GEN_488;
  wire [31:0] _GEN_489;
  wire [31:0] _GEN_490;
  wire [31:0] _GEN_491;
  wire [31:0] _GEN_492;
  wire [31:0] _GEN_493;
  wire [31:0] _GEN_494;
  wire [31:0] _GEN_495;
  wire [31:0] _GEN_496;
  wire [31:0] _GEN_497;
  wire [31:0] _GEN_498;
  wire [31:0] _GEN_499;
  wire [31:0] _GEN_500;
  wire [31:0] _GEN_501;
  wire [31:0] _GEN_502;
  wire [31:0] _GEN_503;
  wire [31:0] _GEN_504;
  wire [31:0] _GEN_505;
  wire [31:0] _GEN_506;
  wire [31:0] _GEN_507;
  wire [31:0] _GEN_508;
  wire [31:0] _GEN_509;
  wire [31:0] _GEN_510;
  wire [31:0] _GEN_511;
  wire [31:0] _GEN_512;
  wire [31:0] _GEN_513;
  wire [31:0] _GEN_514;
  wire [31:0] _GEN_515;
  wire [31:0] _GEN_516;
  wire [31:0] _GEN_517;
  wire [31:0] _GEN_518;
  wire [31:0] _GEN_519;
  wire [31:0] _GEN_520;
  wire [31:0] _GEN_521;
  wire [31:0] _GEN_522;
  wire [31:0] _GEN_523;
  wire [31:0] _GEN_524;
  wire [31:0] _GEN_525;
  wire [31:0] _GEN_526;
  wire [31:0] _GEN_527;
  wire [31:0] _GEN_528;
  wire [31:0] _GEN_529;
  wire [31:0] _GEN_530;
  wire [31:0] _GEN_531;
  wire [31:0] _GEN_532;
  wire [31:0] _GEN_533;
  wire [31:0] _GEN_534;
  wire [31:0] _GEN_535;
  wire [31:0] _GEN_536;
  wire [31:0] _GEN_537;
  wire [31:0] _GEN_538;
  wire [31:0] _GEN_539;
  wire [31:0] _GEN_540;
  wire [31:0] _GEN_541;
  wire [31:0] _GEN_542;
  wire [31:0] _GEN_543;
  wire [31:0] _GEN_544;
  wire [31:0] _GEN_545;
  wire [31:0] _GEN_546;
  wire [31:0] _GEN_547;
  wire [31:0] _GEN_548;
  wire [31:0] _GEN_549;
  wire [31:0] _GEN_550;
  wire [31:0] _GEN_551;
  wire [31:0] _GEN_552;
  wire [31:0] _GEN_553;
  wire [31:0] _GEN_554;
  wire [31:0] _GEN_555;
  wire [31:0] _GEN_556;
  wire [31:0] _GEN_557;
  wire [31:0] _GEN_558;
  wire [31:0] _GEN_559;
  wire [31:0] _GEN_560;
  wire [31:0] _GEN_561;
  wire [31:0] _GEN_562;
  wire [31:0] _GEN_563;
  wire [31:0] _GEN_564;
  wire [31:0] _GEN_565;
  wire [31:0] _GEN_566;
  wire [31:0] _GEN_567;
  wire [31:0] _GEN_568;
  wire [31:0] _GEN_569;
  wire [31:0] _GEN_570;
  wire [31:0] _GEN_571;
  wire [31:0] _GEN_572;
  wire [31:0] _GEN_573;
  wire [31:0] _GEN_574;
  wire [31:0] _GEN_575;
  wire [31:0] _GEN_576;
  wire [31:0] _GEN_577;
  wire [31:0] _GEN_578;
  wire [31:0] _GEN_579;
  wire [31:0] _GEN_580;
  wire [31:0] _GEN_581;
  wire [31:0] _GEN_582;
  wire [31:0] _GEN_583;
  wire [31:0] _GEN_584;
  wire [31:0] _GEN_585;
  wire [31:0] _GEN_586;
  wire [31:0] _GEN_587;
  wire [31:0] _GEN_588;
  wire [31:0] _GEN_589;
  wire [31:0] _GEN_590;
  wire [31:0] _GEN_591;
  wire [31:0] _GEN_592;
  wire [31:0] _GEN_593;
  wire [31:0] _GEN_594;
  wire [31:0] _GEN_595;
  wire [31:0] _GEN_596;
  wire [31:0] _GEN_597;
  wire [31:0] _GEN_598;
  wire [31:0] _GEN_599;
  wire [31:0] _GEN_600;
  wire [31:0] _GEN_601;
  wire [31:0] _GEN_602;
  wire [31:0] _GEN_603;
  wire [31:0] _GEN_604;
  wire [31:0] _GEN_605;
  wire [31:0] _GEN_606;
  wire [31:0] _GEN_607;
  wire [31:0] _GEN_608;
  wire [31:0] _GEN_609;
  wire [31:0] _GEN_610;
  wire [31:0] _GEN_611;
  wire [31:0] _GEN_612;
  wire [31:0] _GEN_613;
  wire [31:0] _GEN_614;
  wire [31:0] _GEN_615;
  wire [31:0] _GEN_616;
  wire [31:0] _GEN_617;
  wire [31:0] _GEN_618;
  wire [31:0] _GEN_619;
  wire [31:0] _GEN_620;
  wire [31:0] _GEN_621;
  wire [31:0] _GEN_622;
  wire [31:0] _GEN_623;
  wire [31:0] _GEN_624;
  wire [31:0] _GEN_625;
  wire [31:0] _GEN_626;
  wire [31:0] _GEN_627;
  wire [31:0] _GEN_628;
  wire [31:0] _GEN_629;
  wire [31:0] _GEN_630;
  wire [31:0] _GEN_631;
  wire [31:0] _GEN_632;
  wire [31:0] _GEN_633;
  wire [31:0] _GEN_634;
  wire [31:0] _GEN_635;
  wire [31:0] _GEN_636;
  wire [31:0] _GEN_637;
  wire [31:0] _GEN_638;
  wire [31:0] _GEN_639;
  wire [31:0] _GEN_640;
  wire [31:0] _GEN_641;
  wire [31:0] _GEN_642;
  wire [31:0] _GEN_643;
  wire [31:0] _GEN_644;
  wire [31:0] _GEN_645;
  wire [31:0] _GEN_646;
  wire [31:0] _GEN_647;
  wire [31:0] _GEN_648;
  wire [31:0] _GEN_649;
  wire [31:0] _GEN_650;
  wire [31:0] _GEN_651;
  wire [31:0] _GEN_652;
  wire [31:0] _GEN_653;
  wire [31:0] _GEN_654;
  wire [31:0] _GEN_655;
  wire [31:0] _GEN_656;
  wire [31:0] _GEN_657;
  wire [31:0] _GEN_658;
  wire [31:0] _GEN_659;
  wire [31:0] _GEN_660;
  wire [31:0] _GEN_661;
  wire [31:0] _GEN_662;
  wire [31:0] _GEN_663;
  wire [31:0] _GEN_664;
  wire [31:0] _GEN_665;
  wire [31:0] _GEN_666;
  wire [31:0] _GEN_667;
  wire [31:0] _GEN_668;
  wire [31:0] _GEN_669;
  wire [31:0] _GEN_670;
  wire [31:0] _GEN_671;
  wire [31:0] _GEN_672;
  wire [31:0] _GEN_673;
  wire [31:0] _GEN_674;
  wire [31:0] _GEN_675;
  wire [31:0] _GEN_676;
  wire [31:0] _GEN_677;
  wire [31:0] _GEN_678;
  wire [31:0] _GEN_679;
  wire [31:0] _GEN_680;
  wire [31:0] _GEN_681;
  wire [31:0] _GEN_682;
  wire [31:0] _GEN_683;
  wire [31:0] _GEN_684;
  wire [31:0] _GEN_685;
  wire [31:0] _GEN_686;
  wire [31:0] _GEN_687;
  wire [31:0] _GEN_688;
  wire [31:0] _GEN_689;
  wire [31:0] _GEN_690;
  wire [31:0] _GEN_691;
  wire [31:0] _GEN_692;
  wire [31:0] _GEN_693;
  wire [31:0] _GEN_694;
  wire [31:0] _GEN_695;
  wire [31:0] _GEN_696;
  wire [31:0] _GEN_697;
  wire [31:0] _GEN_698;
  wire [31:0] _GEN_699;
  wire [31:0] _GEN_700;
  wire [31:0] _GEN_701;
  wire [31:0] _GEN_702;
  wire [31:0] _GEN_703;
  wire [31:0] _GEN_704;
  wire [31:0] _GEN_705;
  wire [31:0] _GEN_706;
  wire [31:0] _GEN_707;
  wire [31:0] _GEN_708;
  wire [31:0] _GEN_709;
  wire [31:0] _GEN_710;
  wire [31:0] _GEN_711;
  wire [31:0] _GEN_712;
  wire [31:0] _GEN_713;
  wire [31:0] _GEN_714;
  wire [31:0] _GEN_715;
  wire [31:0] _GEN_716;
  wire [31:0] _GEN_717;
  wire [31:0] _GEN_718;
  wire [31:0] _GEN_719;
  wire [31:0] _GEN_720;
  wire [31:0] _GEN_721;
  wire [31:0] _GEN_722;
  wire [31:0] _GEN_723;
  wire [31:0] _GEN_724;
  wire [31:0] _GEN_725;
  wire [31:0] _GEN_726;
  wire [31:0] _GEN_727;
  wire [31:0] _GEN_728;
  wire [31:0] _GEN_729;
  wire [31:0] _GEN_730;
  wire [31:0] _GEN_731;
  wire [31:0] _GEN_732;
  wire [31:0] _GEN_733;
  wire [31:0] _GEN_734;
  wire [31:0] _GEN_735;
  wire [31:0] _GEN_736;
  wire [31:0] _GEN_737;
  wire [31:0] _GEN_738;
  wire [31:0] _GEN_739;
  wire [31:0] _GEN_740;
  wire [31:0] _GEN_741;
  wire [31:0] _GEN_742;
  wire [31:0] _GEN_743;
  wire [31:0] _GEN_744;
  wire [31:0] _GEN_745;
  wire [31:0] _GEN_746;
  wire [31:0] _GEN_747;
  wire [31:0] _GEN_748;
  wire [31:0] _GEN_749;
  wire [31:0] _GEN_750;
  wire [31:0] _GEN_751;
  wire [31:0] _GEN_752;
  wire [31:0] _GEN_753;
  wire [31:0] _GEN_754;
  wire [31:0] _GEN_755;
  wire [31:0] _GEN_756;
  wire [31:0] _GEN_757;
  wire [31:0] _GEN_758;
  wire [31:0] _GEN_759;
  wire [31:0] _GEN_760;
  wire [31:0] _GEN_761;
  wire [31:0] _GEN_762;
  wire [31:0] _GEN_763;
  wire [31:0] _GEN_764;
  wire [31:0] _GEN_765;
  wire [31:0] _GEN_766;
  wire [31:0] _GEN_767;
  wire [31:0] _GEN_768;
  wire [31:0] _GEN_769;
  wire [31:0] _GEN_770;
  wire [31:0] _GEN_771;
  wire [31:0] _GEN_772;
  wire [31:0] _GEN_773;
  wire [31:0] _GEN_774;
  wire [31:0] _GEN_775;
  wire [31:0] _GEN_776;
  wire [31:0] _GEN_777;
  wire [31:0] _GEN_778;
  wire [31:0] _GEN_779;
  wire [31:0] _GEN_780;
  wire [31:0] _GEN_781;
  wire [31:0] _GEN_782;
  wire [31:0] _GEN_783;
  wire [31:0] _GEN_784;
  wire [31:0] _GEN_785;
  wire [31:0] _GEN_786;
  wire [31:0] _GEN_787;
  wire [31:0] _GEN_788;
  wire [31:0] _GEN_789;
  wire [31:0] _GEN_790;
  wire [31:0] _GEN_791;
  wire [31:0] _GEN_792;
  wire [31:0] _GEN_793;
  wire [31:0] _GEN_794;
  wire [31:0] _GEN_795;
  wire [31:0] _GEN_796;
  wire [31:0] _GEN_797;
  wire [31:0] _GEN_798;
  wire [31:0] _GEN_799;
  wire [31:0] _GEN_800;
  wire [31:0] _GEN_801;
  wire [31:0] _GEN_802;
  wire [31:0] _GEN_803;
  wire [31:0] _GEN_804;
  wire [31:0] _GEN_805;
  wire [31:0] _GEN_806;
  wire [31:0] _GEN_807;
  wire [31:0] _GEN_808;
  wire [31:0] _GEN_809;
  wire [31:0] _GEN_810;
  wire [31:0] _GEN_811;
  wire [31:0] _GEN_812;
  wire [31:0] _GEN_813;
  wire [31:0] _GEN_814;
  wire [31:0] _GEN_815;
  wire [31:0] _GEN_816;
  wire [31:0] _GEN_817;
  wire [31:0] _GEN_818;
  wire [31:0] _GEN_819;
  wire [31:0] _GEN_820;
  wire [31:0] _GEN_821;
  wire [31:0] _GEN_822;
  wire [31:0] _GEN_823;
  wire [31:0] _GEN_824;
  wire [31:0] _GEN_825;
  wire [31:0] _GEN_826;
  wire [31:0] _GEN_827;
  wire [31:0] _GEN_828;
  wire [31:0] _GEN_829;
  wire [31:0] _GEN_830;
  wire [31:0] _GEN_831;
  wire [31:0] _GEN_832;
  wire [31:0] _GEN_833;
  wire [31:0] _GEN_834;
  wire [31:0] _GEN_835;
  wire [31:0] _GEN_836;
  wire [31:0] _GEN_837;
  wire [31:0] _GEN_838;
  wire [31:0] _GEN_839;
  wire [31:0] _GEN_840;
  wire [31:0] _GEN_841;
  wire [31:0] _GEN_842;
  wire [31:0] _GEN_843;
  wire [31:0] _GEN_844;
  wire [31:0] _GEN_845;
  wire [31:0] _GEN_846;
  wire [31:0] _GEN_847;
  wire [31:0] _GEN_848;
  wire [31:0] _GEN_849;
  wire [31:0] _GEN_850;
  wire [31:0] _GEN_851;
  wire [31:0] _GEN_852;
  wire [31:0] _GEN_853;
  wire [31:0] _GEN_854;
  wire [31:0] _GEN_855;
  wire [31:0] _GEN_856;
  wire [31:0] _GEN_857;
  wire [31:0] _GEN_858;
  wire [31:0] _GEN_859;
  wire [31:0] _GEN_860;
  wire [31:0] _GEN_861;
  wire [31:0] _GEN_862;
  wire [31:0] _GEN_863;
  wire [31:0] _GEN_864;
  wire [31:0] _GEN_865;
  wire [31:0] _GEN_866;
  wire [31:0] _GEN_867;
  wire [31:0] _GEN_868;
  wire [31:0] _GEN_869;
  wire [31:0] _GEN_870;
  wire [31:0] _GEN_871;
  wire [31:0] _GEN_872;
  wire [31:0] _GEN_873;
  wire [31:0] _GEN_874;
  wire [31:0] _GEN_875;
  wire [31:0] _GEN_876;
  wire [31:0] _GEN_877;
  wire [31:0] _GEN_878;
  wire [31:0] _GEN_879;
  wire [31:0] _GEN_880;
  wire [31:0] _GEN_881;
  wire [31:0] _GEN_882;
  wire [31:0] _GEN_883;
  wire [31:0] _GEN_884;
  wire [31:0] _GEN_885;
  wire [31:0] _GEN_886;
  wire [31:0] _GEN_887;
  wire [31:0] _GEN_888;
  wire [31:0] _GEN_889;
  wire [31:0] _GEN_890;
  wire [31:0] _GEN_891;
  wire [31:0] _GEN_892;
  wire [31:0] _GEN_893;
  wire [31:0] _GEN_894;
  wire [31:0] _GEN_895;
  wire [31:0] _GEN_896;
  wire [31:0] _GEN_897;
  wire [31:0] _GEN_898;
  wire [31:0] _GEN_899;
  wire [31:0] _GEN_900;
  wire [31:0] _GEN_901;
  wire [31:0] _GEN_902;
  wire [31:0] _GEN_903;
  wire [31:0] _GEN_904;
  wire [31:0] _GEN_905;
  wire [31:0] _GEN_906;
  wire [31:0] _GEN_907;
  wire [31:0] _GEN_908;
  wire [31:0] _GEN_909;
  wire [31:0] _GEN_910;
  wire [31:0] _GEN_911;
  wire [31:0] _GEN_912;
  wire [31:0] _GEN_913;
  wire [31:0] _GEN_914;
  wire [31:0] _GEN_915;
  wire [31:0] _GEN_916;
  wire [31:0] _GEN_917;
  wire [31:0] _GEN_918;
  wire [31:0] _GEN_919;
  wire [31:0] _GEN_920;
  wire [31:0] _GEN_921;
  wire [31:0] _GEN_922;
  wire [31:0] _GEN_923;
  wire [31:0] _GEN_924;
  wire [31:0] _GEN_925;
  wire [31:0] _GEN_926;
  wire [31:0] _GEN_927;
  wire [31:0] _GEN_928;
  wire [31:0] _GEN_929;
  wire [31:0] _GEN_930;
  wire [31:0] _GEN_931;
  wire [31:0] _GEN_932;
  wire [31:0] _GEN_933;
  wire [31:0] _GEN_934;
  wire [31:0] _GEN_935;
  wire [31:0] _GEN_936;
  wire [31:0] _GEN_937;
  wire [31:0] _GEN_938;
  wire [31:0] _GEN_939;
  wire [31:0] _GEN_940;
  wire [31:0] _GEN_941;
  wire [31:0] _GEN_942;
  wire [31:0] _GEN_943;
  wire [31:0] _GEN_944;
  wire [31:0] _GEN_945;
  wire [31:0] _GEN_946;
  wire [31:0] _GEN_947;
  wire [31:0] _GEN_948;
  wire [31:0] _GEN_949;
  wire [31:0] _GEN_950;
  wire [31:0] _GEN_951;
  wire [31:0] _GEN_952;
  wire [31:0] _GEN_953;
  wire [31:0] _GEN_954;
  wire [31:0] _GEN_955;
  wire [31:0] _GEN_956;
  wire [31:0] _GEN_957;
  wire [31:0] _GEN_958;
  wire [31:0] _GEN_959;
  wire [31:0] _GEN_960;
  wire [31:0] _GEN_961;
  wire [31:0] _GEN_962;
  wire [31:0] _GEN_963;
  wire [31:0] _GEN_964;
  wire [31:0] _GEN_965;
  wire [31:0] _GEN_966;
  wire [31:0] _GEN_967;
  wire [31:0] _GEN_968;
  wire [31:0] _GEN_969;
  wire [31:0] _GEN_970;
  wire [31:0] _GEN_971;
  wire [31:0] _GEN_972;
  wire [31:0] _GEN_973;
  wire [31:0] _GEN_974;
  wire [31:0] _GEN_975;
  wire [31:0] _GEN_976;
  wire [31:0] _GEN_977;
  wire [31:0] _GEN_978;
  wire [31:0] _GEN_979;
  wire [31:0] _GEN_980;
  wire [31:0] _GEN_981;
  wire [31:0] _GEN_982;
  wire [31:0] _GEN_983;
  wire [31:0] _GEN_984;
  wire [31:0] _GEN_985;
  wire [31:0] _GEN_986;
  wire [31:0] _GEN_987;
  wire [31:0] _GEN_988;
  wire [31:0] _GEN_989;
  wire [31:0] _GEN_990;
  wire [31:0] _GEN_991;
  wire [31:0] _GEN_992;
  wire [31:0] _GEN_993;
  wire [31:0] _GEN_994;
  wire [31:0] _GEN_995;
  wire [31:0] _GEN_996;
  wire [31:0] _GEN_997;
  wire [31:0] _GEN_998;
  wire [31:0] _GEN_999;
  wire [31:0] _GEN_1000;
  wire [31:0] _GEN_1001;
  wire [31:0] _GEN_1002;
  wire [31:0] _GEN_1003;
  wire [31:0] _GEN_1004;
  wire [31:0] _GEN_1005;
  wire [31:0] _GEN_1006;
  wire [31:0] _GEN_1007;
  wire [31:0] _GEN_1008;
  wire [31:0] _GEN_1009;
  wire [31:0] _GEN_1010;
  wire [31:0] _GEN_1011;
  wire [31:0] _GEN_1012;
  wire [31:0] _GEN_1013;
  wire [31:0] _GEN_1014;
  wire [31:0] _GEN_1015;
  wire [31:0] _GEN_1016;
  wire [31:0] _GEN_1017;
  wire [31:0] _GEN_1018;
  wire [31:0] _GEN_1019;
  wire [31:0] _GEN_1020;
  wire [31:0] _GEN_1021;
  wire [31:0] _GEN_1022;
  wire [31:0] _GEN_1023;
  wire [31:0] _GEN_1024;
  wire [31:0] _GEN_1025;
  wire [31:0] _GEN_1026;
  wire [31:0] _GEN_1027;
  wire [31:0] _GEN_1028;
  wire [31:0] _GEN_1029;
  wire [31:0] _GEN_1030;
  wire [31:0] _GEN_1031;
  wire [31:0] _GEN_1032;
  wire [31:0] _GEN_1033;
  wire [31:0] _GEN_1034;
  wire [31:0] _GEN_1035;
  wire [31:0] _GEN_1036;
  wire [31:0] _GEN_1037;
  wire [31:0] _GEN_1038;
  wire [31:0] _GEN_1039;
  wire [31:0] _GEN_1040;
  wire [31:0] _GEN_1041;
  wire [31:0] _GEN_1042;
  wire [31:0] _GEN_1043;
  wire [31:0] _GEN_1044;
  wire [31:0] _GEN_1045;
  wire [31:0] _GEN_1046;
  wire [31:0] _GEN_1047;
  wire [31:0] _GEN_1048;
  wire [31:0] _GEN_1049;
  wire [31:0] _GEN_1050;
  wire [31:0] _GEN_1051;
  wire [31:0] _GEN_1052;
  wire [31:0] _GEN_1053;
  wire [31:0] _GEN_1054;
  wire [31:0] _GEN_1055;
  wire [31:0] _GEN_1056;
  wire [31:0] _GEN_1057;
  wire [31:0] _GEN_1058;
  wire [31:0] _GEN_1059;
  wire [31:0] _GEN_1060;
  wire [31:0] _GEN_1061;
  wire [31:0] _GEN_1062;
  wire [31:0] _GEN_1063;
  wire [31:0] _GEN_1064;
  wire [31:0] _GEN_1065;
  wire [31:0] _GEN_1066;
  wire [31:0] _GEN_1067;
  wire [31:0] _GEN_1068;
  wire [31:0] _GEN_1069;
  wire [31:0] _GEN_1070;
  wire [31:0] _GEN_1071;
  wire [31:0] _GEN_1072;
  wire [31:0] _GEN_1073;
  wire [31:0] _GEN_1074;
  wire [31:0] _GEN_1075;
  wire [31:0] _GEN_1076;
  wire [31:0] _GEN_1077;
  wire [31:0] _GEN_1078;
  wire [31:0] _GEN_1079;
  wire [31:0] _GEN_1080;
  wire [31:0] _GEN_1081;
  wire [31:0] _GEN_1082;
  wire [31:0] _GEN_1083;
  wire [31:0] _GEN_1084;
  wire [31:0] _GEN_1085;
  wire [31:0] _GEN_1086;
  wire [31:0] _GEN_1087;
  wire [31:0] _GEN_1088;
  wire [31:0] _GEN_1089;
  wire [31:0] _GEN_1090;
  wire [31:0] _GEN_1091;
  wire [31:0] _GEN_1092;
  wire [31:0] _GEN_1093;
  wire [31:0] _GEN_1094;
  wire [31:0] _GEN_1095;
  wire [31:0] _GEN_1096;
  wire [31:0] _GEN_1097;
  wire [31:0] _GEN_1098;
  wire [31:0] _GEN_1099;
  wire [31:0] _GEN_1100;
  wire [31:0] _GEN_1101;
  wire [31:0] _GEN_1102;
  wire [31:0] _GEN_1103;
  wire [31:0] _GEN_1104;
  wire [31:0] _GEN_1105;
  wire [31:0] _GEN_1106;
  wire [31:0] _GEN_1107;
  wire [31:0] _GEN_1108;
  wire [31:0] _GEN_1109;
  wire [31:0] _GEN_1110;
  wire [31:0] _GEN_1111;
  wire [31:0] _GEN_1112;
  wire [31:0] _GEN_1113;
  wire [31:0] _GEN_1114;
  wire [31:0] _GEN_1115;
  wire [31:0] _GEN_1116;
  wire [31:0] _GEN_1117;
  wire [31:0] _GEN_1118;
  wire [31:0] _GEN_1119;
  wire [31:0] _GEN_1120;
  wire [31:0] _GEN_1121;
  wire [31:0] _GEN_1122;
  wire [31:0] _GEN_1123;
  wire [31:0] _GEN_1124;
  wire [31:0] _GEN_1125;
  wire [31:0] _GEN_1126;
  wire [31:0] _GEN_1127;
  wire [31:0] _GEN_1128;
  wire [31:0] _GEN_1129;
  wire [31:0] _GEN_1130;
  wire [31:0] _GEN_1131;
  wire [31:0] _GEN_1132;
  wire [31:0] _GEN_1133;
  wire [31:0] _GEN_1134;
  wire [31:0] _GEN_1135;
  wire [31:0] _GEN_1136;
  wire [31:0] _GEN_1137;
  wire [31:0] _GEN_1138;
  wire [31:0] _GEN_1139;
  wire [31:0] _GEN_1140;
  wire [31:0] _GEN_1141;
  wire [31:0] _GEN_1142;
  wire [31:0] _GEN_1143;
  wire [31:0] _GEN_1144;
  wire [31:0] _GEN_1145;
  wire [31:0] _GEN_1146;
  wire [31:0] _GEN_1147;
  wire [31:0] _GEN_1148;
  wire [31:0] _GEN_1149;
  wire [31:0] _GEN_1150;
  wire [31:0] _GEN_1151;
  wire [31:0] _GEN_1152;
  wire [31:0] _GEN_1153;
  wire [31:0] _GEN_1154;
  wire [31:0] _GEN_1155;
  wire [31:0] _GEN_1156;
  wire [31:0] _GEN_1157;
  wire [31:0] _GEN_1158;
  wire [31:0] _GEN_1159;
  wire [31:0] _GEN_1160;
  wire [31:0] _GEN_1161;
  wire [31:0] _GEN_1162;
  wire [31:0] _GEN_1163;
  wire [31:0] _GEN_1164;
  wire [31:0] _GEN_1165;
  wire [31:0] _GEN_1166;
  wire [31:0] _GEN_1167;
  wire [31:0] _GEN_1168;
  wire [31:0] _GEN_1169;
  wire [31:0] _GEN_1170;
  wire [31:0] _GEN_1171;
  wire [31:0] _GEN_1172;
  wire [31:0] _GEN_1173;
  wire [31:0] _GEN_1174;
  wire [31:0] _GEN_1175;
  wire [31:0] _GEN_1176;
  wire [31:0] _GEN_1177;
  wire [31:0] _GEN_1178;
  wire [31:0] _GEN_1179;
  wire [31:0] _GEN_1180;
  wire [31:0] _GEN_1181;
  wire [31:0] _GEN_1182;
  wire [31:0] _GEN_1183;
  wire [31:0] _GEN_1184;
  wire [31:0] _GEN_1185;
  wire [31:0] _GEN_1186;
  wire [31:0] _GEN_1187;
  wire [31:0] _GEN_1188;
  wire [31:0] _GEN_1189;
  wire [31:0] _GEN_1190;
  wire [31:0] _GEN_1191;
  wire [31:0] _GEN_1192;
  wire [31:0] _GEN_1193;
  wire [31:0] _GEN_1194;
  wire [31:0] _GEN_1195;
  wire [31:0] _GEN_1196;
  wire [31:0] _GEN_1197;
  wire [31:0] _GEN_1198;
  wire [31:0] _GEN_1199;
  wire [31:0] _GEN_1200;
  wire [31:0] _GEN_1201;
  wire [31:0] _GEN_1202;
  wire [31:0] _GEN_1203;
  wire [31:0] _GEN_1204;
  wire [31:0] _GEN_1205;
  wire [31:0] _GEN_1206;
  wire [31:0] _GEN_1207;
  wire [31:0] _GEN_1208;
  wire [31:0] _GEN_1209;
  wire [31:0] _GEN_1210;
  wire [31:0] _GEN_1211;
  wire [31:0] _GEN_1212;
  wire [31:0] _GEN_1213;
  wire [31:0] _GEN_1214;
  wire [31:0] _GEN_1215;
  wire [31:0] _GEN_1216;
  wire [31:0] _GEN_1217;
  wire [31:0] _GEN_1218;
  wire [31:0] _GEN_1219;
  wire [31:0] _GEN_1220;
  wire [31:0] _GEN_1221;
  wire [31:0] _GEN_1222;
  wire [31:0] _GEN_1223;
  wire [31:0] _GEN_1224;
  wire [31:0] _GEN_1225;
  wire [31:0] _GEN_1226;
  wire [31:0] _GEN_1227;
  wire [31:0] _GEN_1228;
  wire [31:0] _GEN_1229;
  wire [31:0] _GEN_1230;
  wire [31:0] _GEN_1231;
  wire [31:0] _GEN_1232;
  wire [31:0] _GEN_1233;
  wire [31:0] _GEN_1234;
  wire [31:0] _GEN_1235;
  wire [31:0] _GEN_1236;
  wire [31:0] _GEN_1237;
  wire [31:0] _GEN_1238;
  wire [31:0] _GEN_1239;
  wire [31:0] _GEN_1240;
  wire [31:0] _GEN_1241;
  wire [31:0] _GEN_1242;
  wire [31:0] _GEN_1243;
  wire [31:0] _GEN_1244;
  wire [31:0] _GEN_1245;
  wire [31:0] _GEN_1246;
  wire [31:0] _GEN_1247;
  wire [31:0] _GEN_1248;
  wire [31:0] _GEN_1249;
  wire [31:0] _GEN_1250;
  wire [31:0] _GEN_1251;
  wire [31:0] _GEN_1252;
  wire [31:0] _GEN_1253;
  wire [31:0] _GEN_1254;
  wire [31:0] _GEN_1255;
  wire [31:0] _GEN_1256;
  wire [31:0] _GEN_1257;
  wire [31:0] _GEN_1258;
  wire [31:0] _GEN_1259;
  wire [31:0] _GEN_1260;
  wire [31:0] _GEN_1261;
  wire [31:0] _GEN_1262;
  wire [31:0] _GEN_1263;
  wire [31:0] _GEN_1264;
  wire [31:0] _GEN_1265;
  wire [31:0] _GEN_1266;
  wire [31:0] _GEN_1267;
  wire [31:0] _GEN_1268;
  wire [31:0] _GEN_1269;
  wire [31:0] _GEN_1270;
  wire [31:0] _GEN_1271;
  wire [31:0] _GEN_1272;
  wire [31:0] _GEN_1273;
  wire [31:0] _GEN_1274;
  wire [31:0] _GEN_1275;
  wire [31:0] _GEN_1276;
  wire [31:0] _GEN_1277;
  wire [31:0] _GEN_1278;
  wire [31:0] _GEN_1279;
  wire [31:0] _GEN_1280;
  wire [31:0] _GEN_1281;
  wire [31:0] _GEN_1282;
  wire [31:0] _GEN_1283;
  wire [31:0] _GEN_1284;
  wire [31:0] _GEN_1285;
  wire [31:0] _GEN_1286;
  wire [31:0] _GEN_1287;
  wire [31:0] _GEN_1288;
  wire [31:0] _GEN_1289;
  wire [31:0] _GEN_1290;
  wire [31:0] _GEN_1291;
  wire [31:0] _GEN_1292;
  wire [31:0] _GEN_1293;
  wire [31:0] _GEN_1294;
  wire [31:0] _GEN_1295;
  wire [31:0] _GEN_1296;
  wire [31:0] _GEN_1297;
  wire [31:0] _GEN_1298;
  wire [31:0] _GEN_1299;
  wire [31:0] _GEN_1300;
  wire [31:0] _GEN_1301;
  wire [31:0] _GEN_1302;
  wire [31:0] _GEN_1303;
  wire [31:0] _GEN_1304;
  wire [31:0] _GEN_1305;
  wire [31:0] _GEN_1306;
  wire [31:0] _GEN_1307;
  wire [31:0] _GEN_1308;
  wire [31:0] _GEN_1309;
  wire [31:0] _GEN_1310;
  wire [31:0] _GEN_1311;
  wire [31:0] _GEN_1312;
  wire [31:0] _GEN_1313;
  wire [31:0] _GEN_1314;
  wire [31:0] _GEN_1315;
  wire [31:0] _GEN_1316;
  wire [31:0] _GEN_1317;
  wire [31:0] _GEN_1318;
  wire [31:0] _GEN_1319;
  wire [31:0] _GEN_1320;
  wire [31:0] _GEN_1321;
  wire [31:0] _GEN_1322;
  wire [31:0] _GEN_1323;
  wire [31:0] _GEN_1324;
  wire [31:0] _GEN_1325;
  wire [31:0] _GEN_1326;
  wire [31:0] _GEN_1327;
  wire [31:0] _GEN_1328;
  wire [31:0] _GEN_1329;
  wire [31:0] _GEN_1330;
  wire [31:0] _GEN_1331;
  wire [31:0] _GEN_1332;
  wire [31:0] _GEN_1333;
  wire [31:0] _GEN_1334;
  wire [31:0] _GEN_1335;
  wire [31:0] _GEN_1336;
  wire [31:0] _GEN_1337;
  wire [31:0] _GEN_1338;
  wire [31:0] _GEN_1339;
  wire [31:0] _GEN_1340;
  wire [31:0] _GEN_1341;
  wire [31:0] _GEN_1342;
  wire [31:0] _GEN_1343;
  wire [31:0] _GEN_1344;
  wire [31:0] _GEN_1345;
  wire [31:0] _GEN_1346;
  wire [31:0] _GEN_1347;
  wire [31:0] _GEN_1348;
  wire [31:0] _GEN_1349;
  wire [31:0] _GEN_1350;
  wire [31:0] _GEN_1351;
  wire [31:0] _GEN_1352;
  wire [31:0] _GEN_1353;
  wire [31:0] _GEN_1354;
  wire [31:0] _GEN_1355;
  wire [31:0] _GEN_1356;
  wire [31:0] _GEN_1357;
  wire [31:0] _GEN_1358;
  wire [31:0] _GEN_1359;
  wire [31:0] _GEN_1360;
  wire [31:0] _GEN_1361;
  wire [31:0] _GEN_1362;
  wire [31:0] _GEN_1363;
  wire [31:0] _GEN_1364;
  wire [31:0] _GEN_1365;
  wire [31:0] _GEN_1366;
  wire [31:0] _GEN_1367;
  wire [31:0] _GEN_1368;
  wire [31:0] _GEN_1369;
  wire [31:0] _GEN_1370;
  wire [31:0] _GEN_1371;
  wire [31:0] _GEN_1372;
  wire [31:0] _GEN_1373;
  wire [31:0] _GEN_1374;
  wire [31:0] _GEN_1375;
  wire [31:0] _GEN_1376;
  wire [31:0] _GEN_1377;
  wire [31:0] _GEN_1378;
  wire [31:0] _GEN_1379;
  wire [31:0] _GEN_1380;
  wire [31:0] _GEN_1381;
  wire [31:0] _GEN_1382;
  wire [31:0] _GEN_1383;
  wire [31:0] _GEN_1384;
  wire [31:0] _GEN_1385;
  wire [31:0] _GEN_1386;
  wire [31:0] _GEN_1387;
  wire [31:0] _GEN_1388;
  wire [31:0] _GEN_1389;
  wire [31:0] _GEN_1390;
  wire [31:0] _GEN_1391;
  wire [31:0] _GEN_1392;
  wire [31:0] _GEN_1393;
  wire [31:0] _GEN_1394;
  wire [31:0] _GEN_1395;
  wire [31:0] _GEN_1396;
  wire [31:0] _GEN_1397;
  wire [31:0] _GEN_1398;
  wire [31:0] _GEN_1399;
  wire [31:0] _GEN_1400;
  wire [31:0] _GEN_1401;
  wire [31:0] _GEN_1402;
  wire [31:0] _GEN_1403;
  wire [31:0] _GEN_1404;
  wire [31:0] _GEN_1405;
  wire [31:0] _GEN_1406;
  wire [31:0] _GEN_1407;
  wire [31:0] _GEN_1408;
  wire [31:0] _GEN_1409;
  wire [31:0] _GEN_1410;
  wire [31:0] _GEN_1411;
  wire [31:0] _GEN_1412;
  wire [31:0] _GEN_1413;
  wire [31:0] _GEN_1414;
  wire [31:0] _GEN_1415;
  wire [31:0] _GEN_1416;
  wire [31:0] _GEN_1417;
  wire [31:0] _GEN_1418;
  wire [31:0] _GEN_1419;
  wire [31:0] _GEN_1420;
  wire [31:0] _GEN_1421;
  wire [31:0] _GEN_1422;
  wire [31:0] _GEN_1423;
  wire [31:0] _GEN_1424;
  wire [31:0] _GEN_1425;
  wire [31:0] _GEN_1426;
  wire [31:0] _GEN_1427;
  wire [31:0] _GEN_1428;
  wire [31:0] _GEN_1429;
  wire [31:0] _GEN_1430;
  wire [31:0] _GEN_1431;
  wire [31:0] _GEN_1432;
  wire [31:0] _GEN_1433;
  wire [31:0] _GEN_1434;
  wire [31:0] _GEN_1435;
  wire [31:0] _GEN_1436;
  wire [31:0] _GEN_1437;
  wire [31:0] _GEN_1438;
  wire [31:0] _GEN_1439;
  wire [31:0] _GEN_1440;
  wire [31:0] _GEN_1441;
  wire [31:0] _GEN_1442;
  wire [31:0] _GEN_1443;
  wire [31:0] _GEN_1444;
  wire [31:0] _GEN_1445;
  wire [31:0] _GEN_1446;
  wire [31:0] _GEN_1447;
  wire [31:0] _GEN_1448;
  wire [31:0] _GEN_1449;
  wire [31:0] _GEN_1450;
  wire [31:0] _GEN_1451;
  wire [31:0] _GEN_1452;
  wire [31:0] _GEN_1453;
  wire [31:0] _GEN_1454;
  wire [31:0] _GEN_1455;
  wire [31:0] _GEN_1456;
  wire [31:0] _GEN_1457;
  wire [31:0] _GEN_1458;
  wire [31:0] _GEN_1459;
  wire [31:0] _GEN_1460;
  wire [31:0] _GEN_1461;
  wire [31:0] _GEN_1462;
  wire [31:0] _GEN_1463;
  wire [31:0] _GEN_1464;
  wire [31:0] _GEN_1465;
  wire [31:0] _GEN_1466;
  wire [31:0] _GEN_1467;
  wire [31:0] _GEN_1468;
  wire [31:0] _GEN_1469;
  wire [31:0] _GEN_1470;
  wire [31:0] _GEN_1471;
  wire [31:0] _GEN_1472;
  wire [31:0] _GEN_1473;
  wire [31:0] _GEN_1474;
  wire [31:0] _GEN_1475;
  wire [31:0] _GEN_1476;
  wire [31:0] _GEN_1477;
  wire [31:0] _GEN_1478;
  wire [31:0] _GEN_1479;
  wire [31:0] _GEN_1480;
  wire [31:0] _GEN_1481;
  wire [31:0] _GEN_1482;
  wire [31:0] _GEN_1483;
  wire [31:0] _GEN_1484;
  wire [31:0] _GEN_1485;
  wire [31:0] _GEN_1486;
  wire [31:0] _GEN_1487;
  wire [31:0] _GEN_1488;
  wire [31:0] _GEN_1489;
  wire [31:0] _GEN_1490;
  wire [31:0] _GEN_1491;
  wire [31:0] _GEN_1492;
  wire [31:0] _GEN_1493;
  wire [31:0] _GEN_1494;
  wire [31:0] _GEN_1495;
  wire [31:0] _GEN_1496;
  wire [31:0] _GEN_1497;
  wire [31:0] _GEN_1498;
  wire [31:0] _GEN_1499;
  wire [31:0] _GEN_1500;
  wire [31:0] _GEN_1501;
  wire [31:0] _GEN_1502;
  wire [31:0] _GEN_1503;
  wire [31:0] _GEN_1504;
  wire [31:0] _GEN_1505;
  wire [31:0] _GEN_1506;
  wire [31:0] _GEN_1507;
  wire [31:0] _GEN_1508;
  wire [31:0] _GEN_1509;
  wire [31:0] _GEN_1510;
  wire [31:0] _GEN_1511;
  wire [31:0] _GEN_1512;
  wire [31:0] _GEN_1513;
  wire [31:0] _GEN_1514;
  wire [31:0] _GEN_1515;
  wire [31:0] _GEN_1516;
  wire [31:0] _GEN_1517;
  wire [31:0] _GEN_1518;
  wire [31:0] _GEN_1519;
  wire [31:0] _GEN_1520;
  wire [31:0] _GEN_1521;
  wire [31:0] _GEN_1522;
  wire [31:0] _GEN_1523;
  wire [31:0] _GEN_1524;
  wire [31:0] _GEN_1525;
  wire [31:0] _GEN_1526;
  wire [31:0] _GEN_1527;
  wire [31:0] _GEN_1528;
  wire [31:0] _GEN_1529;
  wire [31:0] _GEN_1530;
  wire [31:0] _GEN_1531;
  wire [31:0] _GEN_1532;
  wire [31:0] _GEN_1533;
  wire [31:0] _GEN_1534;
  wire [31:0] _GEN_1535;
  wire [31:0] _GEN_1536;
  wire [31:0] _GEN_1537;
  wire [31:0] _GEN_1538;
  wire [31:0] _GEN_1539;
  wire [31:0] _GEN_1540;
  wire [31:0] _GEN_1541;
  wire [31:0] _GEN_1542;
  wire [31:0] _GEN_1543;
  wire [31:0] _GEN_1544;
  wire [31:0] _GEN_1545;
  wire [31:0] _GEN_1546;
  wire [31:0] _GEN_1547;
  wire [31:0] _GEN_1548;
  wire [31:0] _GEN_1549;
  wire [31:0] _GEN_1550;
  wire [31:0] _GEN_1551;
  wire [31:0] _GEN_1552;
  wire [31:0] _GEN_1553;
  wire [31:0] _GEN_1554;
  wire [31:0] _GEN_1555;
  wire [31:0] _GEN_1556;
  wire [31:0] _GEN_1557;
  wire [31:0] _GEN_1558;
  wire [31:0] _GEN_1559;
  wire [31:0] _GEN_1560;
  wire [31:0] _GEN_1561;
  wire [31:0] _GEN_1562;
  wire [31:0] _GEN_1563;
  wire [31:0] _GEN_1564;
  wire [31:0] _GEN_1565;
  wire [31:0] _GEN_1566;
  wire [31:0] _GEN_1567;
  wire [31:0] _GEN_1568;
  wire [31:0] _GEN_1569;
  wire [31:0] _GEN_1570;
  wire [31:0] _GEN_1571;
  wire [31:0] _GEN_1572;
  wire [31:0] _GEN_1573;
  wire [31:0] _GEN_1574;
  wire [31:0] _GEN_1575;
  wire [31:0] _GEN_1576;
  wire [31:0] _GEN_1577;
  wire [31:0] _GEN_1578;
  wire [31:0] _GEN_1579;
  wire [31:0] _GEN_1580;
  wire [31:0] _GEN_1581;
  wire [31:0] _GEN_1582;
  wire [31:0] _GEN_1583;
  wire [31:0] _GEN_1584;
  wire [31:0] _GEN_1585;
  wire [31:0] _GEN_1586;
  wire [31:0] _GEN_1587;
  wire [31:0] _GEN_1588;
  wire [31:0] _GEN_1589;
  wire [31:0] _GEN_1590;
  wire [31:0] _GEN_1591;
  wire [31:0] _GEN_1592;
  wire [31:0] _GEN_1593;
  wire [31:0] _GEN_1594;
  wire [31:0] _GEN_1595;
  wire [31:0] _GEN_1596;
  wire [31:0] _GEN_1597;
  wire [31:0] _GEN_1598;
  wire [31:0] _GEN_1599;
  wire [31:0] _GEN_1600;
  wire [31:0] _GEN_1601;
  wire [31:0] _GEN_1602;
  wire [31:0] _GEN_1603;
  wire [31:0] _GEN_1604;
  wire [31:0] _GEN_1605;
  wire [31:0] _GEN_1606;
  wire [31:0] _GEN_1607;
  wire [31:0] _GEN_1608;
  wire [31:0] _GEN_1609;
  wire [31:0] _GEN_1610;
  wire [31:0] _GEN_1611;
  wire [31:0] _GEN_1612;
  wire [31:0] _GEN_1613;
  wire [31:0] _GEN_1614;
  wire [31:0] _GEN_1615;
  wire [31:0] _GEN_1616;
  wire [31:0] _GEN_1617;
  wire [31:0] _GEN_1618;
  wire [31:0] _GEN_1619;
  wire [31:0] _GEN_1620;
  wire [31:0] _GEN_1621;
  wire [31:0] _GEN_1622;
  wire [31:0] _GEN_1623;
  wire [31:0] _GEN_1624;
  wire [31:0] _GEN_1625;
  wire [31:0] _GEN_1626;
  wire [31:0] _GEN_1627;
  wire [31:0] _GEN_1628;
  wire [31:0] _GEN_1629;
  wire [31:0] _GEN_1630;
  wire [31:0] _GEN_1631;
  wire [31:0] _GEN_1632;
  wire [31:0] _GEN_1633;
  wire [31:0] _GEN_1634;
  wire [31:0] _GEN_1635;
  wire [31:0] _GEN_1636;
  wire [31:0] _GEN_1637;
  wire [31:0] _GEN_1638;
  wire [31:0] _GEN_1639;
  wire [31:0] _GEN_1640;
  wire [31:0] _GEN_1641;
  wire [31:0] _GEN_1642;
  wire [31:0] _GEN_1643;
  wire [31:0] _GEN_1644;
  wire [31:0] _GEN_1645;
  wire [31:0] _GEN_1646;
  wire [31:0] _GEN_1647;
  wire [31:0] _GEN_1648;
  wire [31:0] _GEN_1649;
  wire [31:0] _GEN_1650;
  wire [31:0] _GEN_1651;
  wire [31:0] _GEN_1652;
  wire [31:0] _GEN_1653;
  wire [31:0] _GEN_1654;
  wire [31:0] _GEN_1655;
  wire [31:0] _GEN_1656;
  wire [31:0] _GEN_1657;
  wire [31:0] _GEN_1658;
  wire [31:0] _GEN_1659;
  wire [31:0] _GEN_1660;
  wire [31:0] _GEN_1661;
  wire [31:0] _GEN_1662;
  wire [31:0] _GEN_1663;
  wire [31:0] _GEN_1664;
  wire [31:0] _GEN_1665;
  wire [31:0] _GEN_1666;
  wire [31:0] _GEN_1667;
  wire [31:0] _GEN_1668;
  wire [31:0] _GEN_1669;
  wire [31:0] _GEN_1670;
  wire [31:0] _GEN_1671;
  wire [31:0] _GEN_1672;
  wire [31:0] _GEN_1673;
  wire [31:0] _GEN_1674;
  wire [31:0] _GEN_1675;
  wire [31:0] _GEN_1676;
  wire [31:0] _GEN_1677;
  wire [31:0] _GEN_1678;
  wire [31:0] _GEN_1679;
  wire [31:0] _GEN_1680;
  wire [31:0] _GEN_1681;
  wire [31:0] _GEN_1682;
  wire [31:0] _GEN_1683;
  wire [31:0] _GEN_1684;
  wire [31:0] _GEN_1685;
  wire [31:0] _GEN_1686;
  wire [31:0] _GEN_1687;
  wire [31:0] _GEN_1688;
  wire [31:0] _GEN_1689;
  wire [31:0] _GEN_1690;
  wire [31:0] _GEN_1691;
  wire [31:0] _GEN_1692;
  wire [31:0] _GEN_1693;
  wire [31:0] _GEN_1694;
  wire [31:0] _GEN_1695;
  wire [31:0] _GEN_1696;
  wire [31:0] _GEN_1697;
  wire [31:0] _GEN_1698;
  wire [31:0] _GEN_1699;
  wire [31:0] _GEN_1700;
  wire [31:0] _GEN_1701;
  wire [31:0] _GEN_1702;
  wire [31:0] _GEN_1703;
  wire [31:0] _GEN_1704;
  wire [31:0] _GEN_1705;
  wire [31:0] _GEN_1706;
  wire [31:0] _GEN_1707;
  wire [31:0] _GEN_1708;
  wire [31:0] _GEN_1709;
  wire [31:0] _GEN_1710;
  wire [31:0] _GEN_1711;
  wire [31:0] _GEN_1712;
  wire [31:0] _GEN_1713;
  wire [31:0] _GEN_1714;
  wire [31:0] _GEN_1715;
  wire [31:0] _GEN_1716;
  wire [31:0] _GEN_1717;
  wire [31:0] _GEN_1718;
  wire [31:0] _GEN_1719;
  wire [31:0] _GEN_1720;
  wire [31:0] _GEN_1721;
  wire [31:0] _GEN_1722;
  wire [31:0] _GEN_1723;
  wire [31:0] _GEN_1724;
  wire [31:0] _GEN_1725;
  wire [31:0] _GEN_1726;
  wire [31:0] _GEN_1727;
  wire [31:0] _GEN_1728;
  wire [31:0] _GEN_1729;
  wire [31:0] _GEN_1730;
  wire [31:0] _GEN_1731;
  wire [31:0] _GEN_1732;
  wire [31:0] _GEN_1733;
  wire [31:0] _GEN_1734;
  wire [31:0] _GEN_1735;
  wire [31:0] _GEN_1736;
  wire [31:0] _GEN_1737;
  wire [31:0] _GEN_1738;
  wire [31:0] _GEN_1739;
  wire [31:0] _GEN_1740;
  wire [31:0] _GEN_1741;
  wire [31:0] _GEN_1742;
  wire [31:0] _GEN_1743;
  wire [31:0] _GEN_1744;
  wire [31:0] _GEN_1745;
  wire [31:0] _GEN_1746;
  wire [31:0] _GEN_1747;
  wire [31:0] _GEN_1748;
  wire [31:0] _GEN_1749;
  wire [31:0] _GEN_1750;
  wire [31:0] _GEN_1751;
  wire [31:0] _GEN_1752;
  wire [31:0] _GEN_1753;
  wire [31:0] _GEN_1754;
  wire [31:0] _GEN_1755;
  wire [31:0] _GEN_1756;
  wire [31:0] _GEN_1757;
  wire [31:0] _GEN_1758;
  wire [31:0] _GEN_1759;
  wire [31:0] _GEN_1760;
  wire [31:0] _GEN_1761;
  wire [31:0] _GEN_1762;
  wire [31:0] _GEN_1763;
  wire [31:0] _GEN_1764;
  wire [31:0] _GEN_1765;
  wire [31:0] _GEN_1766;
  wire [31:0] _GEN_1767;
  wire [31:0] _GEN_1768;
  wire [31:0] _GEN_1769;
  wire [31:0] _GEN_1770;
  wire [31:0] _GEN_1771;
  wire [31:0] _GEN_1772;
  wire [31:0] _GEN_1773;
  wire [31:0] _GEN_1774;
  wire [31:0] _GEN_1775;
  wire [31:0] _GEN_1776;
  wire [31:0] _GEN_1777;
  wire [31:0] _GEN_1778;
  wire [31:0] _GEN_1779;
  wire [31:0] _GEN_1780;
  wire [31:0] _GEN_1781;
  wire [31:0] _GEN_1782;
  wire [31:0] _GEN_1783;
  wire [31:0] _GEN_1784;
  wire [31:0] _GEN_1785;
  wire [31:0] _GEN_1786;
  wire [31:0] _GEN_1787;
  wire [31:0] _GEN_1788;
  wire [31:0] _GEN_1789;
  wire [31:0] _GEN_1790;
  wire [31:0] _GEN_1791;
  wire [31:0] _GEN_1792;
  wire [31:0] _GEN_1793;
  wire [31:0] _GEN_1794;
  wire [31:0] _GEN_1795;
  wire [31:0] _GEN_1796;
  wire [31:0] _GEN_1797;
  wire [31:0] _GEN_1798;
  wire [31:0] _GEN_1799;
  wire [31:0] _GEN_1800;
  wire [31:0] _GEN_1801;
  wire [31:0] _GEN_1802;
  wire [31:0] _GEN_1803;
  wire [31:0] _GEN_1804;
  wire [31:0] _GEN_1805;
  wire [31:0] _GEN_1806;
  wire [31:0] _GEN_1807;
  wire [31:0] _GEN_1808;
  wire [31:0] _GEN_1809;
  wire [31:0] _GEN_1810;
  wire [31:0] _GEN_1811;
  wire [31:0] _GEN_1812;
  wire [31:0] _GEN_1813;
  wire [31:0] _GEN_1814;
  wire [31:0] _GEN_1815;
  wire [31:0] _GEN_1816;
  wire [31:0] _GEN_1817;
  wire [31:0] _GEN_1818;
  wire [31:0] _GEN_1819;
  wire [31:0] _GEN_1820;
  wire [31:0] _GEN_1821;
  wire [31:0] _GEN_1822;
  wire [31:0] _GEN_1823;
  wire [31:0] _GEN_1824;
  wire [31:0] _GEN_1825;
  wire [31:0] _GEN_1826;
  wire [31:0] _GEN_1827;
  wire [31:0] _GEN_1828;
  wire [31:0] _GEN_1829;
  wire [31:0] _GEN_1830;
  wire [31:0] _GEN_1831;
  wire [31:0] _GEN_1832;
  wire [31:0] _GEN_1833;
  wire [31:0] _GEN_1834;
  wire [31:0] _GEN_1835;
  wire [31:0] _GEN_1836;
  wire [31:0] _GEN_1837;
  wire [31:0] _GEN_1838;
  wire [31:0] _GEN_1839;
  wire [31:0] _GEN_1840;
  wire [31:0] _GEN_1841;
  wire [31:0] _GEN_1842;
  wire [31:0] _GEN_1843;
  wire [31:0] _GEN_1844;
  wire [31:0] _GEN_1845;
  wire [31:0] _GEN_1846;
  wire [31:0] _GEN_1847;
  wire [31:0] _GEN_1848;
  wire [31:0] _GEN_1849;
  wire [31:0] _GEN_1850;
  wire [31:0] _GEN_1851;
  wire [31:0] _GEN_1852;
  wire [31:0] _GEN_1853;
  wire [31:0] _GEN_1854;
  wire [31:0] _GEN_1855;
  wire [31:0] _GEN_1856;
  wire [31:0] _GEN_1857;
  wire [31:0] _GEN_1858;
  wire [31:0] _GEN_1859;
  wire [31:0] _GEN_1860;
  wire [31:0] _GEN_1861;
  wire [31:0] _GEN_1862;
  wire [31:0] _GEN_1863;
  wire [31:0] _GEN_1864;
  wire [31:0] _GEN_1865;
  wire [31:0] _GEN_1866;
  wire [31:0] _GEN_1867;
  wire [31:0] _GEN_1868;
  wire [31:0] _GEN_1869;
  wire [31:0] _GEN_1870;
  wire [31:0] _GEN_1871;
  wire [31:0] _GEN_1872;
  wire [31:0] _GEN_1873;
  wire [31:0] _GEN_1874;
  wire [31:0] _GEN_1875;
  wire [31:0] _GEN_1876;
  wire [31:0] _GEN_1877;
  wire [31:0] _GEN_1878;
  wire [31:0] _GEN_1879;
  wire [31:0] _GEN_1880;
  wire [31:0] _GEN_1881;
  wire [31:0] _GEN_1882;
  wire [31:0] _GEN_1883;
  wire [31:0] _GEN_1884;
  wire [31:0] _GEN_1885;
  wire [31:0] _GEN_1886;
  wire [31:0] _GEN_1887;
  wire [31:0] _GEN_1888;
  wire [31:0] _GEN_1889;
  wire [31:0] _GEN_1890;
  wire [31:0] _GEN_1891;
  wire [31:0] _GEN_1892;
  wire [31:0] _GEN_1893;
  wire [31:0] _GEN_1894;
  wire [31:0] _GEN_1895;
  wire [31:0] _GEN_1896;
  wire [31:0] _GEN_1897;
  wire [31:0] _GEN_1898;
  wire [31:0] _GEN_1899;
  wire [31:0] _GEN_1900;
  wire [31:0] _GEN_1901;
  wire [31:0] _GEN_1902;
  wire [31:0] _GEN_1903;
  wire [31:0] _GEN_1904;
  wire [31:0] _GEN_1905;
  wire [31:0] _GEN_1906;
  wire [31:0] _GEN_1907;
  wire [31:0] _GEN_1908;
  wire [31:0] _GEN_1909;
  wire [31:0] _GEN_1910;
  wire [31:0] _GEN_1911;
  wire [31:0] _GEN_1912;
  wire [31:0] _GEN_1913;
  wire [31:0] _GEN_1914;
  wire [31:0] _GEN_1915;
  wire [31:0] _GEN_1916;
  wire [31:0] _GEN_1917;
  wire [31:0] _GEN_1918;
  wire [31:0] _GEN_1919;
  wire [31:0] _GEN_1920;
  wire [31:0] _GEN_1921;
  wire [31:0] _GEN_1922;
  wire [31:0] _GEN_1923;
  wire [31:0] _GEN_1924;
  wire [31:0] _GEN_1925;
  wire [31:0] _GEN_1926;
  wire [31:0] _GEN_1927;
  wire [31:0] _GEN_1928;
  wire [31:0] _GEN_1929;
  wire [31:0] _GEN_1930;
  wire [31:0] _GEN_1931;
  wire [31:0] _GEN_1932;
  wire [31:0] _GEN_1933;
  wire [31:0] _GEN_1934;
  wire [31:0] _GEN_1935;
  wire [31:0] _GEN_1936;
  wire [31:0] _GEN_1937;
  wire [31:0] _GEN_1938;
  wire [31:0] _GEN_1939;
  wire [31:0] _GEN_1940;
  wire [31:0] _GEN_1941;
  wire [31:0] _GEN_1942;
  wire [31:0] _GEN_1943;
  wire [31:0] _GEN_1944;
  wire [31:0] _GEN_1945;
  wire [31:0] _GEN_1946;
  wire [31:0] _GEN_1947;
  wire [31:0] _GEN_1948;
  wire [31:0] _GEN_1949;
  wire [31:0] _GEN_1950;
  wire [31:0] _GEN_1951;
  wire [31:0] _GEN_1952;
  wire [31:0] _GEN_1953;
  wire [31:0] _GEN_1954;
  wire [31:0] _GEN_1955;
  wire [31:0] _GEN_1956;
  wire [31:0] _GEN_1957;
  wire [31:0] _GEN_1958;
  wire [31:0] _GEN_1959;
  wire [31:0] _GEN_1960;
  wire [31:0] _GEN_1961;
  wire [31:0] _GEN_1962;
  wire [31:0] _GEN_1963;
  wire [31:0] _GEN_1964;
  wire [31:0] _GEN_1965;
  wire [31:0] _GEN_1966;
  wire [31:0] _GEN_1967;
  wire [31:0] _GEN_1968;
  wire [31:0] _GEN_1969;
  wire [31:0] _GEN_1970;
  wire [31:0] _GEN_1971;
  wire [31:0] _GEN_1972;
  wire [31:0] _GEN_1973;
  wire [31:0] _GEN_1974;
  wire [31:0] _GEN_1975;
  wire [31:0] _GEN_1976;
  wire [31:0] _GEN_1977;
  wire [31:0] _GEN_1978;
  wire [31:0] _GEN_1979;
  wire [31:0] _GEN_1980;
  wire [31:0] _GEN_1981;
  wire [31:0] _GEN_1982;
  wire [31:0] _GEN_1983;
  wire [31:0] _GEN_1984;
  wire [31:0] _GEN_1985;
  wire [31:0] _GEN_1986;
  wire [31:0] _GEN_1987;
  wire [31:0] _GEN_1988;
  wire [31:0] _GEN_1989;
  wire [31:0] _GEN_1990;
  wire [31:0] _GEN_1991;
  wire [31:0] _GEN_1992;
  wire [31:0] _GEN_1993;
  wire [31:0] _GEN_1994;
  wire [31:0] _GEN_1995;
  wire [31:0] _GEN_1996;
  wire [31:0] _GEN_1997;
  wire [31:0] _GEN_1998;
  wire [31:0] _GEN_1999;
  wire [31:0] _GEN_2000;
  wire [31:0] _GEN_2001;
  wire [31:0] _GEN_2002;
  wire [31:0] _GEN_2003;
  wire [31:0] _GEN_2004;
  wire [31:0] _GEN_2005;
  wire [31:0] _GEN_2006;
  wire [31:0] _GEN_2007;
  wire [31:0] _GEN_2008;
  wire [31:0] _GEN_2009;
  wire [31:0] _GEN_2010;
  wire [31:0] _GEN_2011;
  wire [31:0] _GEN_2012;
  wire [31:0] _GEN_2013;
  wire [31:0] _GEN_2014;
  wire [31:0] _GEN_2015;
  wire [31:0] _GEN_2016;
  wire [31:0] _GEN_2017;
  wire [31:0] _GEN_2018;
  wire [31:0] _GEN_2019;
  wire [31:0] _GEN_2020;
  wire [31:0] _GEN_2021;
  wire [31:0] _GEN_2022;
  wire [31:0] _GEN_2023;
  wire [31:0] _GEN_2024;
  wire [31:0] _GEN_2025;
  wire [31:0] _GEN_2026;
  wire [31:0] _GEN_2027;
  wire [31:0] _GEN_2028;
  wire [31:0] _GEN_2029;
  wire [31:0] _GEN_2030;
  wire [31:0] _GEN_2031;
  wire [31:0] _GEN_2032;
  wire [31:0] _GEN_2033;
  wire [31:0] _GEN_2034;
  wire [31:0] _GEN_2035;
  wire [31:0] _GEN_2036;
  wire [31:0] _GEN_2037;
  wire [31:0] _GEN_2038;
  wire [31:0] _GEN_2039;
  wire [31:0] _GEN_2040;
  wire [31:0] _GEN_2041;
  wire [31:0] _GEN_2042;
  wire [31:0] _GEN_2043;
  wire [31:0] _GEN_2044;
  wire [31:0] _GEN_2045;
  wire [31:0] _GEN_2046;
  wire [31:0] _GEN_2047;
  wire [31:0] _GEN_2048;
  wire [31:0] _GEN_2049;
  wire [31:0] _GEN_2050;
  wire [31:0] _GEN_2051;
  wire [31:0] _GEN_2052;
  wire [7:0] _T_12324;
  wire [7:0] _GEN_2053;
  wire  _T_12325;
  wire [7:0] _T_12328;
  wire [31:0] _GEN_1;
  wire [7:0] _T_12333;
  wire [7:0] _GEN_4101;
  wire  _T_12334;
  wire [7:0] _T_12337;
  wire [31:0] _GEN_2;
  wire [7:0] _T_12342;
  wire [7:0] _GEN_6149;
  wire  _T_12343;
  wire [7:0] _T_12346;
  wire [31:0] _GEN_3;
  wire [7:0] _T_12351;
  wire [7:0] _GEN_8197;
  wire [15:0] _T_12356;
  wire [23:0] _T_12357;
  wire [31:0] _T_12358;
  wire [31:0] _GEN_4;
  wire [31:0] _GEN_8198;
  wire [31:0] _GEN_8199;
  wire [31:0] _GEN_8200;
  wire [31:0] _GEN_8201;
  wire [31:0] _GEN_8202;
  wire [31:0] _GEN_8203;
  wire [31:0] _GEN_8204;
  wire [31:0] _GEN_8205;
  wire [31:0] _GEN_8206;
  wire [31:0] _GEN_8207;
  wire [31:0] _GEN_8208;
  wire [31:0] _GEN_8209;
  wire [31:0] _GEN_8210;
  wire [31:0] _GEN_8211;
  wire [31:0] _GEN_8212;
  wire [31:0] _GEN_8213;
  wire [31:0] _GEN_8214;
  wire [31:0] _GEN_8215;
  wire [31:0] _GEN_8216;
  wire [31:0] _GEN_8217;
  wire [31:0] _GEN_8218;
  wire [31:0] _GEN_8219;
  wire [31:0] _GEN_8220;
  wire [31:0] _GEN_8221;
  wire [31:0] _GEN_8222;
  wire [31:0] _GEN_8223;
  wire [31:0] _GEN_8224;
  wire [31:0] _GEN_8225;
  wire [31:0] _GEN_8226;
  wire [31:0] _GEN_8227;
  wire [31:0] _GEN_8228;
  wire [31:0] _GEN_8229;
  wire [31:0] _GEN_8230;
  wire [31:0] _GEN_8231;
  wire [31:0] _GEN_8232;
  wire [31:0] _GEN_8233;
  wire [31:0] _GEN_8234;
  wire [31:0] _GEN_8235;
  wire [31:0] _GEN_8236;
  wire [31:0] _GEN_8237;
  wire [31:0] _GEN_8238;
  wire [31:0] _GEN_8239;
  wire [31:0] _GEN_8240;
  wire [31:0] _GEN_8241;
  wire [31:0] _GEN_8242;
  wire [31:0] _GEN_8243;
  wire [31:0] _GEN_8244;
  wire [31:0] _GEN_8245;
  wire [31:0] _GEN_8246;
  wire [31:0] _GEN_8247;
  wire [31:0] _GEN_8248;
  wire [31:0] _GEN_8249;
  wire [31:0] _GEN_8250;
  wire [31:0] _GEN_8251;
  wire [31:0] _GEN_8252;
  wire [31:0] _GEN_8253;
  wire [31:0] _GEN_8254;
  wire [31:0] _GEN_8255;
  wire [31:0] _GEN_8256;
  wire [31:0] _GEN_8257;
  wire [31:0] _GEN_8258;
  wire [31:0] _GEN_8259;
  wire [31:0] _GEN_8260;
  wire [31:0] _GEN_8261;
  wire [31:0] _GEN_8262;
  wire [31:0] _GEN_8263;
  wire [31:0] _GEN_8264;
  wire [31:0] _GEN_8265;
  wire [31:0] _GEN_8266;
  wire [31:0] _GEN_8267;
  wire [31:0] _GEN_8268;
  wire [31:0] _GEN_8269;
  wire [31:0] _GEN_8270;
  wire [31:0] _GEN_8271;
  wire [31:0] _GEN_8272;
  wire [31:0] _GEN_8273;
  wire [31:0] _GEN_8274;
  wire [31:0] _GEN_8275;
  wire [31:0] _GEN_8276;
  wire [31:0] _GEN_8277;
  wire [31:0] _GEN_8278;
  wire [31:0] _GEN_8279;
  wire [31:0] _GEN_8280;
  wire [31:0] _GEN_8281;
  wire [31:0] _GEN_8282;
  wire [31:0] _GEN_8283;
  wire [31:0] _GEN_8284;
  wire [31:0] _GEN_8285;
  wire [31:0] _GEN_8286;
  wire [31:0] _GEN_8287;
  wire [31:0] _GEN_8288;
  wire [31:0] _GEN_8289;
  wire [31:0] _GEN_8290;
  wire [31:0] _GEN_8291;
  wire [31:0] _GEN_8292;
  wire [31:0] _GEN_8293;
  wire [31:0] _GEN_8294;
  wire [31:0] _GEN_8295;
  wire [31:0] _GEN_8296;
  wire [31:0] _GEN_8297;
  wire [31:0] _GEN_8298;
  wire [31:0] _GEN_8299;
  wire [31:0] _GEN_8300;
  wire [31:0] _GEN_8301;
  wire [31:0] _GEN_8302;
  wire [31:0] _GEN_8303;
  wire [31:0] _GEN_8304;
  wire [31:0] _GEN_8305;
  wire [31:0] _GEN_8306;
  wire [31:0] _GEN_8307;
  wire [31:0] _GEN_8308;
  wire [31:0] _GEN_8309;
  wire [31:0] _GEN_8310;
  wire [31:0] _GEN_8311;
  wire [31:0] _GEN_8312;
  wire [31:0] _GEN_8313;
  wire [31:0] _GEN_8314;
  wire [31:0] _GEN_8315;
  wire [31:0] _GEN_8316;
  wire [31:0] _GEN_8317;
  wire [31:0] _GEN_8318;
  wire [31:0] _GEN_8319;
  wire [31:0] _GEN_8320;
  wire [31:0] _GEN_8321;
  wire [31:0] _GEN_8322;
  wire [31:0] _GEN_8323;
  wire [31:0] _GEN_8324;
  wire [31:0] _GEN_8325;
  wire [31:0] _GEN_8326;
  wire [31:0] _GEN_8327;
  wire [31:0] _GEN_8328;
  wire [31:0] _GEN_8329;
  wire [31:0] _GEN_8330;
  wire [31:0] _GEN_8331;
  wire [31:0] _GEN_8332;
  wire [31:0] _GEN_8333;
  wire [31:0] _GEN_8334;
  wire [31:0] _GEN_8335;
  wire [31:0] _GEN_8336;
  wire [31:0] _GEN_8337;
  wire [31:0] _GEN_8338;
  wire [31:0] _GEN_8339;
  wire [31:0] _GEN_8340;
  wire [31:0] _GEN_8341;
  wire [31:0] _GEN_8342;
  wire [31:0] _GEN_8343;
  wire [31:0] _GEN_8344;
  wire [31:0] _GEN_8345;
  wire [31:0] _GEN_8346;
  wire [31:0] _GEN_8347;
  wire [31:0] _GEN_8348;
  wire [31:0] _GEN_8349;
  wire [31:0] _GEN_8350;
  wire [31:0] _GEN_8351;
  wire [31:0] _GEN_8352;
  wire [31:0] _GEN_8353;
  wire [31:0] _GEN_8354;
  wire [31:0] _GEN_8355;
  wire [31:0] _GEN_8356;
  wire [31:0] _GEN_8357;
  wire [31:0] _GEN_8358;
  wire [31:0] _GEN_8359;
  wire [31:0] _GEN_8360;
  wire [31:0] _GEN_8361;
  wire [31:0] _GEN_8362;
  wire [31:0] _GEN_8363;
  wire [31:0] _GEN_8364;
  wire [31:0] _GEN_8365;
  wire [31:0] _GEN_8366;
  wire [31:0] _GEN_8367;
  wire [31:0] _GEN_8368;
  wire [31:0] _GEN_8369;
  wire [31:0] _GEN_8370;
  wire [31:0] _GEN_8371;
  wire [31:0] _GEN_8372;
  wire [31:0] _GEN_8373;
  wire [31:0] _GEN_8374;
  wire [31:0] _GEN_8375;
  wire [31:0] _GEN_8376;
  wire [31:0] _GEN_8377;
  wire [31:0] _GEN_8378;
  wire [31:0] _GEN_8379;
  wire [31:0] _GEN_8380;
  wire [31:0] _GEN_8381;
  wire [31:0] _GEN_8382;
  wire [31:0] _GEN_8383;
  wire [31:0] _GEN_8384;
  wire [31:0] _GEN_8385;
  wire [31:0] _GEN_8386;
  wire [31:0] _GEN_8387;
  wire [31:0] _GEN_8388;
  wire [31:0] _GEN_8389;
  wire [31:0] _GEN_8390;
  wire [31:0] _GEN_8391;
  wire [31:0] _GEN_8392;
  wire [31:0] _GEN_8393;
  wire [31:0] _GEN_8394;
  wire [31:0] _GEN_8395;
  wire [31:0] _GEN_8396;
  wire [31:0] _GEN_8397;
  wire [31:0] _GEN_8398;
  wire [31:0] _GEN_8399;
  wire [31:0] _GEN_8400;
  wire [31:0] _GEN_8401;
  wire [31:0] _GEN_8402;
  wire [31:0] _GEN_8403;
  wire [31:0] _GEN_8404;
  wire [31:0] _GEN_8405;
  wire [31:0] _GEN_8406;
  wire [31:0] _GEN_8407;
  wire [31:0] _GEN_8408;
  wire [31:0] _GEN_8409;
  wire [31:0] _GEN_8410;
  wire [31:0] _GEN_8411;
  wire [31:0] _GEN_8412;
  wire [31:0] _GEN_8413;
  wire [31:0] _GEN_8414;
  wire [31:0] _GEN_8415;
  wire [31:0] _GEN_8416;
  wire [31:0] _GEN_8417;
  wire [31:0] _GEN_8418;
  wire [31:0] _GEN_8419;
  wire [31:0] _GEN_8420;
  wire [31:0] _GEN_8421;
  wire [31:0] _GEN_8422;
  wire [31:0] _GEN_8423;
  wire [31:0] _GEN_8424;
  wire [31:0] _GEN_8425;
  wire [31:0] _GEN_8426;
  wire [31:0] _GEN_8427;
  wire [31:0] _GEN_8428;
  wire [31:0] _GEN_8429;
  wire [31:0] _GEN_8430;
  wire [31:0] _GEN_8431;
  wire [31:0] _GEN_8432;
  wire [31:0] _GEN_8433;
  wire [31:0] _GEN_8434;
  wire [31:0] _GEN_8435;
  wire [31:0] _GEN_8436;
  wire [31:0] _GEN_8437;
  wire [31:0] _GEN_8438;
  wire [31:0] _GEN_8439;
  wire [31:0] _GEN_8440;
  wire [31:0] _GEN_8441;
  wire [31:0] _GEN_8442;
  wire [31:0] _GEN_8443;
  wire [31:0] _GEN_8444;
  wire [31:0] _GEN_8445;
  wire [31:0] _GEN_8446;
  wire [31:0] _GEN_8447;
  wire [31:0] _GEN_8448;
  wire [31:0] _GEN_8449;
  wire [31:0] _GEN_8450;
  wire [31:0] _GEN_8451;
  wire [31:0] _GEN_8452;
  wire [31:0] _GEN_8453;
  wire [31:0] _GEN_8454;
  wire [31:0] _GEN_8455;
  wire [31:0] _GEN_8456;
  wire [31:0] _GEN_8457;
  wire [31:0] _GEN_8458;
  wire [31:0] _GEN_8459;
  wire [31:0] _GEN_8460;
  wire [31:0] _GEN_8461;
  wire [31:0] _GEN_8462;
  wire [31:0] _GEN_8463;
  wire [31:0] _GEN_8464;
  wire [31:0] _GEN_8465;
  wire [31:0] _GEN_8466;
  wire [31:0] _GEN_8467;
  wire [31:0] _GEN_8468;
  wire [31:0] _GEN_8469;
  wire [31:0] _GEN_8470;
  wire [31:0] _GEN_8471;
  wire [31:0] _GEN_8472;
  wire [31:0] _GEN_8473;
  wire [31:0] _GEN_8474;
  wire [31:0] _GEN_8475;
  wire [31:0] _GEN_8476;
  wire [31:0] _GEN_8477;
  wire [31:0] _GEN_8478;
  wire [31:0] _GEN_8479;
  wire [31:0] _GEN_8480;
  wire [31:0] _GEN_8481;
  wire [31:0] _GEN_8482;
  wire [31:0] _GEN_8483;
  wire [31:0] _GEN_8484;
  wire [31:0] _GEN_8485;
  wire [31:0] _GEN_8486;
  wire [31:0] _GEN_8487;
  wire [31:0] _GEN_8488;
  wire [31:0] _GEN_8489;
  wire [31:0] _GEN_8490;
  wire [31:0] _GEN_8491;
  wire [31:0] _GEN_8492;
  wire [31:0] _GEN_8493;
  wire [31:0] _GEN_8494;
  wire [31:0] _GEN_8495;
  wire [31:0] _GEN_8496;
  wire [31:0] _GEN_8497;
  wire [31:0] _GEN_8498;
  wire [31:0] _GEN_8499;
  wire [31:0] _GEN_8500;
  wire [31:0] _GEN_8501;
  wire [31:0] _GEN_8502;
  wire [31:0] _GEN_8503;
  wire [31:0] _GEN_8504;
  wire [31:0] _GEN_8505;
  wire [31:0] _GEN_8506;
  wire [31:0] _GEN_8507;
  wire [31:0] _GEN_8508;
  wire [31:0] _GEN_8509;
  wire [31:0] _GEN_8510;
  wire [31:0] _GEN_8511;
  wire [31:0] _GEN_8512;
  wire [31:0] _GEN_8513;
  wire [31:0] _GEN_8514;
  wire [31:0] _GEN_8515;
  wire [31:0] _GEN_8516;
  wire [31:0] _GEN_8517;
  wire [31:0] _GEN_8518;
  wire [31:0] _GEN_8519;
  wire [31:0] _GEN_8520;
  wire [31:0] _GEN_8521;
  wire [31:0] _GEN_8522;
  wire [31:0] _GEN_8523;
  wire [31:0] _GEN_8524;
  wire [31:0] _GEN_8525;
  wire [31:0] _GEN_8526;
  wire [31:0] _GEN_8527;
  wire [31:0] _GEN_8528;
  wire [31:0] _GEN_8529;
  wire [31:0] _GEN_8530;
  wire [31:0] _GEN_8531;
  wire [31:0] _GEN_8532;
  wire [31:0] _GEN_8533;
  wire [31:0] _GEN_8534;
  wire [31:0] _GEN_8535;
  wire [31:0] _GEN_8536;
  wire [31:0] _GEN_8537;
  wire [31:0] _GEN_8538;
  wire [31:0] _GEN_8539;
  wire [31:0] _GEN_8540;
  wire [31:0] _GEN_8541;
  wire [31:0] _GEN_8542;
  wire [31:0] _GEN_8543;
  wire [31:0] _GEN_8544;
  wire [31:0] _GEN_8545;
  wire [31:0] _GEN_8546;
  wire [31:0] _GEN_8547;
  wire [31:0] _GEN_8548;
  wire [31:0] _GEN_8549;
  wire [31:0] _GEN_8550;
  wire [31:0] _GEN_8551;
  wire [31:0] _GEN_8552;
  wire [31:0] _GEN_8553;
  wire [31:0] _GEN_8554;
  wire [31:0] _GEN_8555;
  wire [31:0] _GEN_8556;
  wire [31:0] _GEN_8557;
  wire [31:0] _GEN_8558;
  wire [31:0] _GEN_8559;
  wire [31:0] _GEN_8560;
  wire [31:0] _GEN_8561;
  wire [31:0] _GEN_8562;
  wire [31:0] _GEN_8563;
  wire [31:0] _GEN_8564;
  wire [31:0] _GEN_8565;
  wire [31:0] _GEN_8566;
  wire [31:0] _GEN_8567;
  wire [31:0] _GEN_8568;
  wire [31:0] _GEN_8569;
  wire [31:0] _GEN_8570;
  wire [31:0] _GEN_8571;
  wire [31:0] _GEN_8572;
  wire [31:0] _GEN_8573;
  wire [31:0] _GEN_8574;
  wire [31:0] _GEN_8575;
  wire [31:0] _GEN_8576;
  wire [31:0] _GEN_8577;
  wire [31:0] _GEN_8578;
  wire [31:0] _GEN_8579;
  wire [31:0] _GEN_8580;
  wire [31:0] _GEN_8581;
  wire [31:0] _GEN_8582;
  wire [31:0] _GEN_8583;
  wire [31:0] _GEN_8584;
  wire [31:0] _GEN_8585;
  wire [31:0] _GEN_8586;
  wire [31:0] _GEN_8587;
  wire [31:0] _GEN_8588;
  wire [31:0] _GEN_8589;
  wire [31:0] _GEN_8590;
  wire [31:0] _GEN_8591;
  wire [31:0] _GEN_8592;
  wire [31:0] _GEN_8593;
  wire [31:0] _GEN_8594;
  wire [31:0] _GEN_8595;
  wire [31:0] _GEN_8596;
  wire [31:0] _GEN_8597;
  wire [31:0] _GEN_8598;
  wire [31:0] _GEN_8599;
  wire [31:0] _GEN_8600;
  wire [31:0] _GEN_8601;
  wire [31:0] _GEN_8602;
  wire [31:0] _GEN_8603;
  wire [31:0] _GEN_8604;
  wire [31:0] _GEN_8605;
  wire [31:0] _GEN_8606;
  wire [31:0] _GEN_8607;
  wire [31:0] _GEN_8608;
  wire [31:0] _GEN_8609;
  wire [31:0] _GEN_8610;
  wire [31:0] _GEN_8611;
  wire [31:0] _GEN_8612;
  wire [31:0] _GEN_8613;
  wire [31:0] _GEN_8614;
  wire [31:0] _GEN_8615;
  wire [31:0] _GEN_8616;
  wire [31:0] _GEN_8617;
  wire [31:0] _GEN_8618;
  wire [31:0] _GEN_8619;
  wire [31:0] _GEN_8620;
  wire [31:0] _GEN_8621;
  wire [31:0] _GEN_8622;
  wire [31:0] _GEN_8623;
  wire [31:0] _GEN_8624;
  wire [31:0] _GEN_8625;
  wire [31:0] _GEN_8626;
  wire [31:0] _GEN_8627;
  wire [31:0] _GEN_8628;
  wire [31:0] _GEN_8629;
  wire [31:0] _GEN_8630;
  wire [31:0] _GEN_8631;
  wire [31:0] _GEN_8632;
  wire [31:0] _GEN_8633;
  wire [31:0] _GEN_8634;
  wire [31:0] _GEN_8635;
  wire [31:0] _GEN_8636;
  wire [31:0] _GEN_8637;
  wire [31:0] _GEN_8638;
  wire [31:0] _GEN_8639;
  wire [31:0] _GEN_8640;
  wire [31:0] _GEN_8641;
  wire [31:0] _GEN_8642;
  wire [31:0] _GEN_8643;
  wire [31:0] _GEN_8644;
  wire [31:0] _GEN_8645;
  wire [31:0] _GEN_8646;
  wire [31:0] _GEN_8647;
  wire [31:0] _GEN_8648;
  wire [31:0] _GEN_8649;
  wire [31:0] _GEN_8650;
  wire [31:0] _GEN_8651;
  wire [31:0] _GEN_8652;
  wire [31:0] _GEN_8653;
  wire [31:0] _GEN_8654;
  wire [31:0] _GEN_8655;
  wire [31:0] _GEN_8656;
  wire [31:0] _GEN_8657;
  wire [31:0] _GEN_8658;
  wire [31:0] _GEN_8659;
  wire [31:0] _GEN_8660;
  wire [31:0] _GEN_8661;
  wire [31:0] _GEN_8662;
  wire [31:0] _GEN_8663;
  wire [31:0] _GEN_8664;
  wire [31:0] _GEN_8665;
  wire [31:0] _GEN_8666;
  wire [31:0] _GEN_8667;
  wire [31:0] _GEN_8668;
  wire [31:0] _GEN_8669;
  wire [31:0] _GEN_8670;
  wire [31:0] _GEN_8671;
  wire [31:0] _GEN_8672;
  wire [31:0] _GEN_8673;
  wire [31:0] _GEN_8674;
  wire [31:0] _GEN_8675;
  wire [31:0] _GEN_8676;
  wire [31:0] _GEN_8677;
  wire [31:0] _GEN_8678;
  wire [31:0] _GEN_8679;
  wire [31:0] _GEN_8680;
  wire [31:0] _GEN_8681;
  wire [31:0] _GEN_8682;
  wire [31:0] _GEN_8683;
  wire [31:0] _GEN_8684;
  wire [31:0] _GEN_8685;
  wire [31:0] _GEN_8686;
  wire [31:0] _GEN_8687;
  wire [31:0] _GEN_8688;
  wire [31:0] _GEN_8689;
  wire [31:0] _GEN_8690;
  wire [31:0] _GEN_8691;
  wire [31:0] _GEN_8692;
  wire [31:0] _GEN_8693;
  wire [31:0] _GEN_8694;
  wire [31:0] _GEN_8695;
  wire [31:0] _GEN_8696;
  wire [31:0] _GEN_8697;
  wire [31:0] _GEN_8698;
  wire [31:0] _GEN_8699;
  wire [31:0] _GEN_8700;
  wire [31:0] _GEN_8701;
  wire [31:0] _GEN_8702;
  wire [31:0] _GEN_8703;
  wire [31:0] _GEN_8704;
  wire [31:0] _GEN_8705;
  wire [31:0] _GEN_8706;
  wire [31:0] _GEN_8707;
  wire [31:0] _GEN_8708;
  wire [31:0] _GEN_8709;
  wire [31:0] _GEN_8710;
  wire [31:0] _GEN_8711;
  wire [31:0] _GEN_8712;
  wire [31:0] _GEN_8713;
  wire [31:0] _GEN_8714;
  wire [31:0] _GEN_8715;
  wire [31:0] _GEN_8716;
  wire [31:0] _GEN_8717;
  wire [31:0] _GEN_8718;
  wire [31:0] _GEN_8719;
  wire [31:0] _GEN_8720;
  wire [31:0] _GEN_8721;
  wire [31:0] _GEN_8722;
  wire [31:0] _GEN_8723;
  wire [31:0] _GEN_8724;
  wire [31:0] _GEN_8725;
  wire [31:0] _GEN_8726;
  wire [31:0] _GEN_8727;
  wire [31:0] _GEN_8728;
  wire [31:0] _GEN_8729;
  wire [31:0] _GEN_8730;
  wire [31:0] _GEN_8731;
  wire [31:0] _GEN_8732;
  wire [31:0] _GEN_8733;
  wire [31:0] _GEN_8734;
  wire [31:0] _GEN_8735;
  wire [31:0] _GEN_8736;
  wire [31:0] _GEN_8737;
  wire [31:0] _GEN_8738;
  wire [31:0] _GEN_8739;
  wire [31:0] _GEN_8740;
  wire [31:0] _GEN_8741;
  wire [31:0] _GEN_8742;
  wire [31:0] _GEN_8743;
  wire [31:0] _GEN_8744;
  wire [31:0] _GEN_8745;
  wire [31:0] _GEN_8746;
  wire [31:0] _GEN_8747;
  wire [31:0] _GEN_8748;
  wire [31:0] _GEN_8749;
  wire [31:0] _GEN_8750;
  wire [31:0] _GEN_8751;
  wire [31:0] _GEN_8752;
  wire [31:0] _GEN_8753;
  wire [31:0] _GEN_8754;
  wire [31:0] _GEN_8755;
  wire [31:0] _GEN_8756;
  wire [31:0] _GEN_8757;
  wire [31:0] _GEN_8758;
  wire [31:0] _GEN_8759;
  wire [31:0] _GEN_8760;
  wire [31:0] _GEN_8761;
  wire [31:0] _GEN_8762;
  wire [31:0] _GEN_8763;
  wire [31:0] _GEN_8764;
  wire [31:0] _GEN_8765;
  wire [31:0] _GEN_8766;
  wire [31:0] _GEN_8767;
  wire [31:0] _GEN_8768;
  wire [31:0] _GEN_8769;
  wire [31:0] _GEN_8770;
  wire [31:0] _GEN_8771;
  wire [31:0] _GEN_8772;
  wire [31:0] _GEN_8773;
  wire [31:0] _GEN_8774;
  wire [31:0] _GEN_8775;
  wire [31:0] _GEN_8776;
  wire [31:0] _GEN_8777;
  wire [31:0] _GEN_8778;
  wire [31:0] _GEN_8779;
  wire [31:0] _GEN_8780;
  wire [31:0] _GEN_8781;
  wire [31:0] _GEN_8782;
  wire [31:0] _GEN_8783;
  wire [31:0] _GEN_8784;
  wire [31:0] _GEN_8785;
  wire [31:0] _GEN_8786;
  wire [31:0] _GEN_8787;
  wire [31:0] _GEN_8788;
  wire [31:0] _GEN_8789;
  wire [31:0] _GEN_8790;
  wire [31:0] _GEN_8791;
  wire [31:0] _GEN_8792;
  wire [31:0] _GEN_8793;
  wire [31:0] _GEN_8794;
  wire [31:0] _GEN_8795;
  wire [31:0] _GEN_8796;
  wire [31:0] _GEN_8797;
  wire [31:0] _GEN_8798;
  wire [31:0] _GEN_8799;
  wire [31:0] _GEN_8800;
  wire [31:0] _GEN_8801;
  wire [31:0] _GEN_8802;
  wire [31:0] _GEN_8803;
  wire [31:0] _GEN_8804;
  wire [31:0] _GEN_8805;
  wire [31:0] _GEN_8806;
  wire [31:0] _GEN_8807;
  wire [31:0] _GEN_8808;
  wire [31:0] _GEN_8809;
  wire [31:0] _GEN_8810;
  wire [31:0] _GEN_8811;
  wire [31:0] _GEN_8812;
  wire [31:0] _GEN_8813;
  wire [31:0] _GEN_8814;
  wire [31:0] _GEN_8815;
  wire [31:0] _GEN_8816;
  wire [31:0] _GEN_8817;
  wire [31:0] _GEN_8818;
  wire [31:0] _GEN_8819;
  wire [31:0] _GEN_8820;
  wire [31:0] _GEN_8821;
  wire [31:0] _GEN_8822;
  wire [31:0] _GEN_8823;
  wire [31:0] _GEN_8824;
  wire [31:0] _GEN_8825;
  wire [31:0] _GEN_8826;
  wire [31:0] _GEN_8827;
  wire [31:0] _GEN_8828;
  wire [31:0] _GEN_8829;
  wire [31:0] _GEN_8830;
  wire [31:0] _GEN_8831;
  wire [31:0] _GEN_8832;
  wire [31:0] _GEN_8833;
  wire [31:0] _GEN_8834;
  wire [31:0] _GEN_8835;
  wire [31:0] _GEN_8836;
  wire [31:0] _GEN_8837;
  wire [31:0] _GEN_8838;
  wire [31:0] _GEN_8839;
  wire [31:0] _GEN_8840;
  wire [31:0] _GEN_8841;
  wire [31:0] _GEN_8842;
  wire [31:0] _GEN_8843;
  wire [31:0] _GEN_8844;
  wire [31:0] _GEN_8845;
  wire [31:0] _GEN_8846;
  wire [31:0] _GEN_8847;
  wire [31:0] _GEN_8848;
  wire [31:0] _GEN_8849;
  wire [31:0] _GEN_8850;
  wire [31:0] _GEN_8851;
  wire [31:0] _GEN_8852;
  wire [31:0] _GEN_8853;
  wire [31:0] _GEN_8854;
  wire [31:0] _GEN_8855;
  wire [31:0] _GEN_8856;
  wire [31:0] _GEN_8857;
  wire [31:0] _GEN_8858;
  wire [31:0] _GEN_8859;
  wire [31:0] _GEN_8860;
  wire [31:0] _GEN_8861;
  wire [31:0] _GEN_8862;
  wire [31:0] _GEN_8863;
  wire [31:0] _GEN_8864;
  wire [31:0] _GEN_8865;
  wire [31:0] _GEN_8866;
  wire [31:0] _GEN_8867;
  wire [31:0] _GEN_8868;
  wire [31:0] _GEN_8869;
  wire [31:0] _GEN_8870;
  wire [31:0] _GEN_8871;
  wire [31:0] _GEN_8872;
  wire [31:0] _GEN_8873;
  wire [31:0] _GEN_8874;
  wire [31:0] _GEN_8875;
  wire [31:0] _GEN_8876;
  wire [31:0] _GEN_8877;
  wire [31:0] _GEN_8878;
  wire [31:0] _GEN_8879;
  wire [31:0] _GEN_8880;
  wire [31:0] _GEN_8881;
  wire [31:0] _GEN_8882;
  wire [31:0] _GEN_8883;
  wire [31:0] _GEN_8884;
  wire [31:0] _GEN_8885;
  wire [31:0] _GEN_8886;
  wire [31:0] _GEN_8887;
  wire [31:0] _GEN_8888;
  wire [31:0] _GEN_8889;
  wire [31:0] _GEN_8890;
  wire [31:0] _GEN_8891;
  wire [31:0] _GEN_8892;
  wire [31:0] _GEN_8893;
  wire [31:0] _GEN_8894;
  wire [31:0] _GEN_8895;
  wire [31:0] _GEN_8896;
  wire [31:0] _GEN_8897;
  wire [31:0] _GEN_8898;
  wire [31:0] _GEN_8899;
  wire [31:0] _GEN_8900;
  wire [31:0] _GEN_8901;
  wire [31:0] _GEN_8902;
  wire [31:0] _GEN_8903;
  wire [31:0] _GEN_8904;
  wire [31:0] _GEN_8905;
  wire [31:0] _GEN_8906;
  wire [31:0] _GEN_8907;
  wire [31:0] _GEN_8908;
  wire [31:0] _GEN_8909;
  wire [31:0] _GEN_8910;
  wire [31:0] _GEN_8911;
  wire [31:0] _GEN_8912;
  wire [31:0] _GEN_8913;
  wire [31:0] _GEN_8914;
  wire [31:0] _GEN_8915;
  wire [31:0] _GEN_8916;
  wire [31:0] _GEN_8917;
  wire [31:0] _GEN_8918;
  wire [31:0] _GEN_8919;
  wire [31:0] _GEN_8920;
  wire [31:0] _GEN_8921;
  wire [31:0] _GEN_8922;
  wire [31:0] _GEN_8923;
  wire [31:0] _GEN_8924;
  wire [31:0] _GEN_8925;
  wire [31:0] _GEN_8926;
  wire [31:0] _GEN_8927;
  wire [31:0] _GEN_8928;
  wire [31:0] _GEN_8929;
  wire [31:0] _GEN_8930;
  wire [31:0] _GEN_8931;
  wire [31:0] _GEN_8932;
  wire [31:0] _GEN_8933;
  wire [31:0] _GEN_8934;
  wire [31:0] _GEN_8935;
  wire [31:0] _GEN_8936;
  wire [31:0] _GEN_8937;
  wire [31:0] _GEN_8938;
  wire [31:0] _GEN_8939;
  wire [31:0] _GEN_8940;
  wire [31:0] _GEN_8941;
  wire [31:0] _GEN_8942;
  wire [31:0] _GEN_8943;
  wire [31:0] _GEN_8944;
  wire [31:0] _GEN_8945;
  wire [31:0] _GEN_8946;
  wire [31:0] _GEN_8947;
  wire [31:0] _GEN_8948;
  wire [31:0] _GEN_8949;
  wire [31:0] _GEN_8950;
  wire [31:0] _GEN_8951;
  wire [31:0] _GEN_8952;
  wire [31:0] _GEN_8953;
  wire [31:0] _GEN_8954;
  wire [31:0] _GEN_8955;
  wire [31:0] _GEN_8956;
  wire [31:0] _GEN_8957;
  wire [31:0] _GEN_8958;
  wire [31:0] _GEN_8959;
  wire [31:0] _GEN_8960;
  wire [31:0] _GEN_8961;
  wire [31:0] _GEN_8962;
  wire [31:0] _GEN_8963;
  wire [31:0] _GEN_8964;
  wire [31:0] _GEN_8965;
  wire [31:0] _GEN_8966;
  wire [31:0] _GEN_8967;
  wire [31:0] _GEN_8968;
  wire [31:0] _GEN_8969;
  wire [31:0] _GEN_8970;
  wire [31:0] _GEN_8971;
  wire [31:0] _GEN_8972;
  wire [31:0] _GEN_8973;
  wire [31:0] _GEN_8974;
  wire [31:0] _GEN_8975;
  wire [31:0] _GEN_8976;
  wire [31:0] _GEN_8977;
  wire [31:0] _GEN_8978;
  wire [31:0] _GEN_8979;
  wire [31:0] _GEN_8980;
  wire [31:0] _GEN_8981;
  wire [31:0] _GEN_8982;
  wire [31:0] _GEN_8983;
  wire [31:0] _GEN_8984;
  wire [31:0] _GEN_8985;
  wire [31:0] _GEN_8986;
  wire [31:0] _GEN_8987;
  wire [31:0] _GEN_8988;
  wire [31:0] _GEN_8989;
  wire [31:0] _GEN_8990;
  wire [31:0] _GEN_8991;
  wire [31:0] _GEN_8992;
  wire [31:0] _GEN_8993;
  wire [31:0] _GEN_8994;
  wire [31:0] _GEN_8995;
  wire [31:0] _GEN_8996;
  wire [31:0] _GEN_8997;
  wire [31:0] _GEN_8998;
  wire [31:0] _GEN_8999;
  wire [31:0] _GEN_9000;
  wire [31:0] _GEN_9001;
  wire [31:0] _GEN_9002;
  wire [31:0] _GEN_9003;
  wire [31:0] _GEN_9004;
  wire [31:0] _GEN_9005;
  wire [31:0] _GEN_9006;
  wire [31:0] _GEN_9007;
  wire [31:0] _GEN_9008;
  wire [31:0] _GEN_9009;
  wire [31:0] _GEN_9010;
  wire [31:0] _GEN_9011;
  wire [31:0] _GEN_9012;
  wire [31:0] _GEN_9013;
  wire [31:0] _GEN_9014;
  wire [31:0] _GEN_9015;
  wire [31:0] _GEN_9016;
  wire [31:0] _GEN_9017;
  wire [31:0] _GEN_9018;
  wire [31:0] _GEN_9019;
  wire [31:0] _GEN_9020;
  wire [31:0] _GEN_9021;
  wire [31:0] _GEN_9022;
  wire [31:0] _GEN_9023;
  wire [31:0] _GEN_9024;
  wire [31:0] _GEN_9025;
  wire [31:0] _GEN_9026;
  wire [31:0] _GEN_9027;
  wire [31:0] _GEN_9028;
  wire [31:0] _GEN_9029;
  wire [31:0] _GEN_9030;
  wire [31:0] _GEN_9031;
  wire [31:0] _GEN_9032;
  wire [31:0] _GEN_9033;
  wire [31:0] _GEN_9034;
  wire [31:0] _GEN_9035;
  wire [31:0] _GEN_9036;
  wire [31:0] _GEN_9037;
  wire [31:0] _GEN_9038;
  wire [31:0] _GEN_9039;
  wire [31:0] _GEN_9040;
  wire [31:0] _GEN_9041;
  wire [31:0] _GEN_9042;
  wire [31:0] _GEN_9043;
  wire [31:0] _GEN_9044;
  wire [31:0] _GEN_9045;
  wire [31:0] _GEN_9046;
  wire [31:0] _GEN_9047;
  wire [31:0] _GEN_9048;
  wire [31:0] _GEN_9049;
  wire [31:0] _GEN_9050;
  wire [31:0] _GEN_9051;
  wire [31:0] _GEN_9052;
  wire [31:0] _GEN_9053;
  wire [31:0] _GEN_9054;
  wire [31:0] _GEN_9055;
  wire [31:0] _GEN_9056;
  wire [31:0] _GEN_9057;
  wire [31:0] _GEN_9058;
  wire [31:0] _GEN_9059;
  wire [31:0] _GEN_9060;
  wire [31:0] _GEN_9061;
  wire [31:0] _GEN_9062;
  wire [31:0] _GEN_9063;
  wire [31:0] _GEN_9064;
  wire [31:0] _GEN_9065;
  wire [31:0] _GEN_9066;
  wire [31:0] _GEN_9067;
  wire [31:0] _GEN_9068;
  wire [31:0] _GEN_9069;
  wire [31:0] _GEN_9070;
  wire [31:0] _GEN_9071;
  wire [31:0] _GEN_9072;
  wire [31:0] _GEN_9073;
  wire [31:0] _GEN_9074;
  wire [31:0] _GEN_9075;
  wire [31:0] _GEN_9076;
  wire [31:0] _GEN_9077;
  wire [31:0] _GEN_9078;
  wire [31:0] _GEN_9079;
  wire [31:0] _GEN_9080;
  wire [31:0] _GEN_9081;
  wire [31:0] _GEN_9082;
  wire [31:0] _GEN_9083;
  wire [31:0] _GEN_9084;
  wire [31:0] _GEN_9085;
  wire [31:0] _GEN_9086;
  wire [31:0] _GEN_9087;
  wire [31:0] _GEN_9088;
  wire [31:0] _GEN_9089;
  wire [31:0] _GEN_9090;
  wire [31:0] _GEN_9091;
  wire [31:0] _GEN_9092;
  wire [31:0] _GEN_9093;
  wire [31:0] _GEN_9094;
  wire [31:0] _GEN_9095;
  wire [31:0] _GEN_9096;
  wire [31:0] _GEN_9097;
  wire [31:0] _GEN_9098;
  wire [31:0] _GEN_9099;
  wire [31:0] _GEN_9100;
  wire [31:0] _GEN_9101;
  wire [31:0] _GEN_9102;
  wire [31:0] _GEN_9103;
  wire [31:0] _GEN_9104;
  wire [31:0] _GEN_9105;
  wire [31:0] _GEN_9106;
  wire [31:0] _GEN_9107;
  wire [31:0] _GEN_9108;
  wire [31:0] _GEN_9109;
  wire [31:0] _GEN_9110;
  wire [31:0] _GEN_9111;
  wire [31:0] _GEN_9112;
  wire [31:0] _GEN_9113;
  wire [31:0] _GEN_9114;
  wire [31:0] _GEN_9115;
  wire [31:0] _GEN_9116;
  wire [31:0] _GEN_9117;
  wire [31:0] _GEN_9118;
  wire [31:0] _GEN_9119;
  wire [31:0] _GEN_9120;
  wire [31:0] _GEN_9121;
  wire [31:0] _GEN_9122;
  wire [31:0] _GEN_9123;
  wire [31:0] _GEN_9124;
  wire [31:0] _GEN_9125;
  wire [31:0] _GEN_9126;
  wire [31:0] _GEN_9127;
  wire [31:0] _GEN_9128;
  wire [31:0] _GEN_9129;
  wire [31:0] _GEN_9130;
  wire [31:0] _GEN_9131;
  wire [31:0] _GEN_9132;
  wire [31:0] _GEN_9133;
  wire [31:0] _GEN_9134;
  wire [31:0] _GEN_9135;
  wire [31:0] _GEN_9136;
  wire [31:0] _GEN_9137;
  wire [31:0] _GEN_9138;
  wire [31:0] _GEN_9139;
  wire [31:0] _GEN_9140;
  wire [31:0] _GEN_9141;
  wire [31:0] _GEN_9142;
  wire [31:0] _GEN_9143;
  wire [31:0] _GEN_9144;
  wire [31:0] _GEN_9145;
  wire [31:0] _GEN_9146;
  wire [31:0] _GEN_9147;
  wire [31:0] _GEN_9148;
  wire [31:0] _GEN_9149;
  wire [31:0] _GEN_9150;
  wire [31:0] _GEN_9151;
  wire [31:0] _GEN_9152;
  wire [31:0] _GEN_9153;
  wire [31:0] _GEN_9154;
  wire [31:0] _GEN_9155;
  wire [31:0] _GEN_9156;
  wire [31:0] _GEN_9157;
  wire [31:0] _GEN_9158;
  wire [31:0] _GEN_9159;
  wire [31:0] _GEN_9160;
  wire [31:0] _GEN_9161;
  wire [31:0] _GEN_9162;
  wire [31:0] _GEN_9163;
  wire [31:0] _GEN_9164;
  wire [31:0] _GEN_9165;
  wire [31:0] _GEN_9166;
  wire [31:0] _GEN_9167;
  wire [31:0] _GEN_9168;
  wire [31:0] _GEN_9169;
  wire [31:0] _GEN_9170;
  wire [31:0] _GEN_9171;
  wire [31:0] _GEN_9172;
  wire [31:0] _GEN_9173;
  wire [31:0] _GEN_9174;
  wire [31:0] _GEN_9175;
  wire [31:0] _GEN_9176;
  wire [31:0] _GEN_9177;
  wire [31:0] _GEN_9178;
  wire [31:0] _GEN_9179;
  wire [31:0] _GEN_9180;
  wire [31:0] _GEN_9181;
  wire [31:0] _GEN_9182;
  wire [31:0] _GEN_9183;
  wire [31:0] _GEN_9184;
  wire [31:0] _GEN_9185;
  wire [31:0] _GEN_9186;
  wire [31:0] _GEN_9187;
  wire [31:0] _GEN_9188;
  wire [31:0] _GEN_9189;
  wire [31:0] _GEN_9190;
  wire [31:0] _GEN_9191;
  wire [31:0] _GEN_9192;
  wire [31:0] _GEN_9193;
  wire [31:0] _GEN_9194;
  wire [31:0] _GEN_9195;
  wire [31:0] _GEN_9196;
  wire [31:0] _GEN_9197;
  wire [31:0] _GEN_9198;
  wire [31:0] _GEN_9199;
  wire [31:0] _GEN_9200;
  wire [31:0] _GEN_9201;
  wire [31:0] _GEN_9202;
  wire [31:0] _GEN_9203;
  wire [31:0] _GEN_9204;
  wire [31:0] _GEN_9205;
  wire [31:0] _GEN_9206;
  wire [31:0] _GEN_9207;
  wire [31:0] _GEN_9208;
  wire [31:0] _GEN_9209;
  wire [31:0] _GEN_9210;
  wire [31:0] _GEN_9211;
  wire [31:0] _GEN_9212;
  wire [31:0] _GEN_9213;
  wire [31:0] _GEN_9214;
  wire [31:0] _GEN_9215;
  wire [31:0] _GEN_9216;
  wire [31:0] _GEN_9217;
  wire [31:0] _GEN_9218;
  wire [31:0] _GEN_9219;
  wire [31:0] _GEN_9220;
  wire [31:0] _GEN_9221;
  wire [31:0] _GEN_9222;
  wire [31:0] _GEN_9223;
  wire [31:0] _GEN_9224;
  wire [31:0] _GEN_9225;
  wire [31:0] _GEN_9226;
  wire [31:0] _GEN_9227;
  wire [31:0] _GEN_9228;
  wire [31:0] _GEN_9229;
  wire [31:0] _GEN_9230;
  wire [31:0] _GEN_9231;
  wire [31:0] _GEN_9232;
  wire [31:0] _GEN_9233;
  wire [31:0] _GEN_9234;
  wire [31:0] _GEN_9235;
  wire [31:0] _GEN_9236;
  wire [31:0] _GEN_9237;
  wire [31:0] _GEN_9238;
  wire [31:0] _GEN_9239;
  wire [31:0] _GEN_9240;
  wire [31:0] _GEN_9241;
  wire [31:0] _GEN_9242;
  wire [31:0] _GEN_9243;
  wire [31:0] _GEN_9244;
  wire [31:0] _GEN_9245;
  wire [31:0] _GEN_9246;
  wire [31:0] _GEN_9247;
  wire [31:0] _GEN_9248;
  wire [31:0] _GEN_9249;
  wire [31:0] _GEN_9250;
  wire [31:0] _GEN_9251;
  wire [31:0] _GEN_9252;
  wire [31:0] _GEN_9253;
  wire [31:0] _GEN_9254;
  wire [31:0] _GEN_9255;
  wire [31:0] _GEN_9256;
  wire [31:0] _GEN_9257;
  wire [31:0] _GEN_9258;
  wire [31:0] _GEN_9259;
  wire [31:0] _GEN_9260;
  wire [31:0] _GEN_9261;
  wire [31:0] _GEN_9262;
  wire [31:0] _GEN_9263;
  wire [31:0] _GEN_9264;
  wire [31:0] _GEN_9265;
  wire [31:0] _GEN_9266;
  wire [31:0] _GEN_9267;
  wire [31:0] _GEN_9268;
  wire [31:0] _GEN_9269;
  wire [31:0] _GEN_9270;
  wire [31:0] _GEN_9271;
  wire [31:0] _GEN_9272;
  wire [31:0] _GEN_9273;
  wire [31:0] _GEN_9274;
  wire [31:0] _GEN_9275;
  wire [31:0] _GEN_9276;
  wire [31:0] _GEN_9277;
  wire [31:0] _GEN_9278;
  wire [31:0] _GEN_9279;
  wire [31:0] _GEN_9280;
  wire [31:0] _GEN_9281;
  wire [31:0] _GEN_9282;
  wire [31:0] _GEN_9283;
  wire [31:0] _GEN_9284;
  wire [31:0] _GEN_9285;
  wire [31:0] _GEN_9286;
  wire [31:0] _GEN_9287;
  wire [31:0] _GEN_9288;
  wire [31:0] _GEN_9289;
  wire [31:0] _GEN_9290;
  wire [31:0] _GEN_9291;
  wire [31:0] _GEN_9292;
  wire [31:0] _GEN_9293;
  wire [31:0] _GEN_9294;
  wire [31:0] _GEN_9295;
  wire [31:0] _GEN_9296;
  wire [31:0] _GEN_9297;
  wire [31:0] _GEN_9298;
  wire [31:0] _GEN_9299;
  wire [31:0] _GEN_9300;
  wire [31:0] _GEN_9301;
  wire [31:0] _GEN_9302;
  wire [31:0] _GEN_9303;
  wire [31:0] _GEN_9304;
  wire [31:0] _GEN_9305;
  wire [31:0] _GEN_9306;
  wire [31:0] _GEN_9307;
  wire [31:0] _GEN_9308;
  wire [31:0] _GEN_9309;
  wire [31:0] _GEN_9310;
  wire [31:0] _GEN_9311;
  wire [31:0] _GEN_9312;
  wire [31:0] _GEN_9313;
  wire [31:0] _GEN_9314;
  wire [31:0] _GEN_9315;
  wire [31:0] _GEN_9316;
  wire [31:0] _GEN_9317;
  wire [31:0] _GEN_9318;
  wire [31:0] _GEN_9319;
  wire [31:0] _GEN_9320;
  wire [31:0] _GEN_9321;
  wire [31:0] _GEN_9322;
  wire [31:0] _GEN_9323;
  wire [31:0] _GEN_9324;
  wire [31:0] _GEN_9325;
  wire [31:0] _GEN_9326;
  wire [31:0] _GEN_9327;
  wire [31:0] _GEN_9328;
  wire [31:0] _GEN_9329;
  wire [31:0] _GEN_9330;
  wire [31:0] _GEN_9331;
  wire [31:0] _GEN_9332;
  wire [31:0] _GEN_9333;
  wire [31:0] _GEN_9334;
  wire [31:0] _GEN_9335;
  wire [31:0] _GEN_9336;
  wire [31:0] _GEN_9337;
  wire [31:0] _GEN_9338;
  wire [31:0] _GEN_9339;
  wire [31:0] _GEN_9340;
  wire [31:0] _GEN_9341;
  wire [31:0] _GEN_9342;
  wire [31:0] _GEN_9343;
  wire [31:0] _GEN_9344;
  wire [31:0] _GEN_9345;
  wire [31:0] _GEN_9346;
  wire [31:0] _GEN_9347;
  wire [31:0] _GEN_9348;
  wire [31:0] _GEN_9349;
  wire [31:0] _GEN_9350;
  wire [31:0] _GEN_9351;
  wire [31:0] _GEN_9352;
  wire [31:0] _GEN_9353;
  wire [31:0] _GEN_9354;
  wire [31:0] _GEN_9355;
  wire [31:0] _GEN_9356;
  wire [31:0] _GEN_9357;
  wire [31:0] _GEN_9358;
  wire [31:0] _GEN_9359;
  wire [31:0] _GEN_9360;
  wire [31:0] _GEN_9361;
  wire [31:0] _GEN_9362;
  wire [31:0] _GEN_9363;
  wire [31:0] _GEN_9364;
  wire [31:0] _GEN_9365;
  wire [31:0] _GEN_9366;
  wire [31:0] _GEN_9367;
  wire [31:0] _GEN_9368;
  wire [31:0] _GEN_9369;
  wire [31:0] _GEN_9370;
  wire [31:0] _GEN_9371;
  wire [31:0] _GEN_9372;
  wire [31:0] _GEN_9373;
  wire [31:0] _GEN_9374;
  wire [31:0] _GEN_9375;
  wire [31:0] _GEN_9376;
  wire [31:0] _GEN_9377;
  wire [31:0] _GEN_9378;
  wire [31:0] _GEN_9379;
  wire [31:0] _GEN_9380;
  wire [31:0] _GEN_9381;
  wire [31:0] _GEN_9382;
  wire [31:0] _GEN_9383;
  wire [31:0] _GEN_9384;
  wire [31:0] _GEN_9385;
  wire [31:0] _GEN_9386;
  wire [31:0] _GEN_9387;
  wire [31:0] _GEN_9388;
  wire [31:0] _GEN_9389;
  wire [31:0] _GEN_9390;
  wire [31:0] _GEN_9391;
  wire [31:0] _GEN_9392;
  wire [31:0] _GEN_9393;
  wire [31:0] _GEN_9394;
  wire [31:0] _GEN_9395;
  wire [31:0] _GEN_9396;
  wire [31:0] _GEN_9397;
  wire [31:0] _GEN_9398;
  wire [31:0] _GEN_9399;
  wire [31:0] _GEN_9400;
  wire [31:0] _GEN_9401;
  wire [31:0] _GEN_9402;
  wire [31:0] _GEN_9403;
  wire [31:0] _GEN_9404;
  wire [31:0] _GEN_9405;
  wire [31:0] _GEN_9406;
  wire [31:0] _GEN_9407;
  wire [31:0] _GEN_9408;
  wire [31:0] _GEN_9409;
  wire [31:0] _GEN_9410;
  wire [31:0] _GEN_9411;
  wire [31:0] _GEN_9412;
  wire [31:0] _GEN_9413;
  wire [31:0] _GEN_9414;
  wire [31:0] _GEN_9415;
  wire [31:0] _GEN_9416;
  wire [31:0] _GEN_9417;
  wire [31:0] _GEN_9418;
  wire [31:0] _GEN_9419;
  wire [31:0] _GEN_9420;
  wire [31:0] _GEN_9421;
  wire [31:0] _GEN_9422;
  wire [31:0] _GEN_9423;
  wire [31:0] _GEN_9424;
  wire [31:0] _GEN_9425;
  wire [31:0] _GEN_9426;
  wire [31:0] _GEN_9427;
  wire [31:0] _GEN_9428;
  wire [31:0] _GEN_9429;
  wire [31:0] _GEN_9430;
  wire [31:0] _GEN_9431;
  wire [31:0] _GEN_9432;
  wire [31:0] _GEN_9433;
  wire [31:0] _GEN_9434;
  wire [31:0] _GEN_9435;
  wire [31:0] _GEN_9436;
  wire [31:0] _GEN_9437;
  wire [31:0] _GEN_9438;
  wire [31:0] _GEN_9439;
  wire [31:0] _GEN_9440;
  wire [31:0] _GEN_9441;
  wire [31:0] _GEN_9442;
  wire [31:0] _GEN_9443;
  wire [31:0] _GEN_9444;
  wire [31:0] _GEN_9445;
  wire [31:0] _GEN_9446;
  wire [31:0] _GEN_9447;
  wire [31:0] _GEN_9448;
  wire [31:0] _GEN_9449;
  wire [31:0] _GEN_9450;
  wire [31:0] _GEN_9451;
  wire [31:0] _GEN_9452;
  wire [31:0] _GEN_9453;
  wire [31:0] _GEN_9454;
  wire [31:0] _GEN_9455;
  wire [31:0] _GEN_9456;
  wire [31:0] _GEN_9457;
  wire [31:0] _GEN_9458;
  wire [31:0] _GEN_9459;
  wire [31:0] _GEN_9460;
  wire [31:0] _GEN_9461;
  wire [31:0] _GEN_9462;
  wire [31:0] _GEN_9463;
  wire [31:0] _GEN_9464;
  wire [31:0] _GEN_9465;
  wire [31:0] _GEN_9466;
  wire [31:0] _GEN_9467;
  wire [31:0] _GEN_9468;
  wire [31:0] _GEN_9469;
  wire [31:0] _GEN_9470;
  wire [31:0] _GEN_9471;
  wire [31:0] _GEN_9472;
  wire [31:0] _GEN_9473;
  wire [31:0] _GEN_9474;
  wire [31:0] _GEN_9475;
  wire [31:0] _GEN_9476;
  wire [31:0] _GEN_9477;
  wire [31:0] _GEN_9478;
  wire [31:0] _GEN_9479;
  wire [31:0] _GEN_9480;
  wire [31:0] _GEN_9481;
  wire [31:0] _GEN_9482;
  wire [31:0] _GEN_9483;
  wire [31:0] _GEN_9484;
  wire [31:0] _GEN_9485;
  wire [31:0] _GEN_9486;
  wire [31:0] _GEN_9487;
  wire [31:0] _GEN_9488;
  wire [31:0] _GEN_9489;
  wire [31:0] _GEN_9490;
  wire [31:0] _GEN_9491;
  wire [31:0] _GEN_9492;
  wire [31:0] _GEN_9493;
  wire [31:0] _GEN_9494;
  wire [31:0] _GEN_9495;
  wire [31:0] _GEN_9496;
  wire [31:0] _GEN_9497;
  wire [31:0] _GEN_9498;
  wire [31:0] _GEN_9499;
  wire [31:0] _GEN_9500;
  wire [31:0] _GEN_9501;
  wire [31:0] _GEN_9502;
  wire [31:0] _GEN_9503;
  wire [31:0] _GEN_9504;
  wire [31:0] _GEN_9505;
  wire [31:0] _GEN_9506;
  wire [31:0] _GEN_9507;
  wire [31:0] _GEN_9508;
  wire [31:0] _GEN_9509;
  wire [31:0] _GEN_9510;
  wire [31:0] _GEN_9511;
  wire [31:0] _GEN_9512;
  wire [31:0] _GEN_9513;
  wire [31:0] _GEN_9514;
  wire [31:0] _GEN_9515;
  wire [31:0] _GEN_9516;
  wire [31:0] _GEN_9517;
  wire [31:0] _GEN_9518;
  wire [31:0] _GEN_9519;
  wire [31:0] _GEN_9520;
  wire [31:0] _GEN_9521;
  wire [31:0] _GEN_9522;
  wire [31:0] _GEN_9523;
  wire [31:0] _GEN_9524;
  wire [31:0] _GEN_9525;
  wire [31:0] _GEN_9526;
  wire [31:0] _GEN_9527;
  wire [31:0] _GEN_9528;
  wire [31:0] _GEN_9529;
  wire [31:0] _GEN_9530;
  wire [31:0] _GEN_9531;
  wire [31:0] _GEN_9532;
  wire [31:0] _GEN_9533;
  wire [31:0] _GEN_9534;
  wire [31:0] _GEN_9535;
  wire [31:0] _GEN_9536;
  wire [31:0] _GEN_9537;
  wire [31:0] _GEN_9538;
  wire [31:0] _GEN_9539;
  wire [31:0] _GEN_9540;
  wire [31:0] _GEN_9541;
  wire [31:0] _GEN_9542;
  wire [31:0] _GEN_9543;
  wire [31:0] _GEN_9544;
  wire [31:0] _GEN_9545;
  wire [31:0] _GEN_9546;
  wire [31:0] _GEN_9547;
  wire [31:0] _GEN_9548;
  wire [31:0] _GEN_9549;
  wire [31:0] _GEN_9550;
  wire [31:0] _GEN_9551;
  wire [31:0] _GEN_9552;
  wire [31:0] _GEN_9553;
  wire [31:0] _GEN_9554;
  wire [31:0] _GEN_9555;
  wire [31:0] _GEN_9556;
  wire [31:0] _GEN_9557;
  wire [31:0] _GEN_9558;
  wire [31:0] _GEN_9559;
  wire [31:0] _GEN_9560;
  wire [31:0] _GEN_9561;
  wire [31:0] _GEN_9562;
  wire [31:0] _GEN_9563;
  wire [31:0] _GEN_9564;
  wire [31:0] _GEN_9565;
  wire [31:0] _GEN_9566;
  wire [31:0] _GEN_9567;
  wire [31:0] _GEN_9568;
  wire [31:0] _GEN_9569;
  wire [31:0] _GEN_9570;
  wire [31:0] _GEN_9571;
  wire [31:0] _GEN_9572;
  wire [31:0] _GEN_9573;
  wire [31:0] _GEN_9574;
  wire [31:0] _GEN_9575;
  wire [31:0] _GEN_9576;
  wire [31:0] _GEN_9577;
  wire [31:0] _GEN_9578;
  wire [31:0] _GEN_9579;
  wire [31:0] _GEN_9580;
  wire [31:0] _GEN_9581;
  wire [31:0] _GEN_9582;
  wire [31:0] _GEN_9583;
  wire [31:0] _GEN_9584;
  wire [31:0] _GEN_9585;
  wire [31:0] _GEN_9586;
  wire [31:0] _GEN_9587;
  wire [31:0] _GEN_9588;
  wire [31:0] _GEN_9589;
  wire [31:0] _GEN_9590;
  wire [31:0] _GEN_9591;
  wire [31:0] _GEN_9592;
  wire [31:0] _GEN_9593;
  wire [31:0] _GEN_9594;
  wire [31:0] _GEN_9595;
  wire [31:0] _GEN_9596;
  wire [31:0] _GEN_9597;
  wire [31:0] _GEN_9598;
  wire [31:0] _GEN_9599;
  wire [31:0] _GEN_9600;
  wire [31:0] _GEN_9601;
  wire [31:0] _GEN_9602;
  wire [31:0] _GEN_9603;
  wire [31:0] _GEN_9604;
  wire [31:0] _GEN_9605;
  wire [31:0] _GEN_9606;
  wire [31:0] _GEN_9607;
  wire [31:0] _GEN_9608;
  wire [31:0] _GEN_9609;
  wire [31:0] _GEN_9610;
  wire [31:0] _GEN_9611;
  wire [31:0] _GEN_9612;
  wire [31:0] _GEN_9613;
  wire [31:0] _GEN_9614;
  wire [31:0] _GEN_9615;
  wire [31:0] _GEN_9616;
  wire [31:0] _GEN_9617;
  wire [31:0] _GEN_9618;
  wire [31:0] _GEN_9619;
  wire [31:0] _GEN_9620;
  wire [31:0] _GEN_9621;
  wire [31:0] _GEN_9622;
  wire [31:0] _GEN_9623;
  wire [31:0] _GEN_9624;
  wire [31:0] _GEN_9625;
  wire [31:0] _GEN_9626;
  wire [31:0] _GEN_9627;
  wire [31:0] _GEN_9628;
  wire [31:0] _GEN_9629;
  wire [31:0] _GEN_9630;
  wire [31:0] _GEN_9631;
  wire [31:0] _GEN_9632;
  wire [31:0] _GEN_9633;
  wire [31:0] _GEN_9634;
  wire [31:0] _GEN_9635;
  wire [31:0] _GEN_9636;
  wire [31:0] _GEN_9637;
  wire [31:0] _GEN_9638;
  wire [31:0] _GEN_9639;
  wire [31:0] _GEN_9640;
  wire [31:0] _GEN_9641;
  wire [31:0] _GEN_9642;
  wire [31:0] _GEN_9643;
  wire [31:0] _GEN_9644;
  wire [31:0] _GEN_9645;
  wire [31:0] _GEN_9646;
  wire [31:0] _GEN_9647;
  wire [31:0] _GEN_9648;
  wire [31:0] _GEN_9649;
  wire [31:0] _GEN_9650;
  wire [31:0] _GEN_9651;
  wire [31:0] _GEN_9652;
  wire [31:0] _GEN_9653;
  wire [31:0] _GEN_9654;
  wire [31:0] _GEN_9655;
  wire [31:0] _GEN_9656;
  wire [31:0] _GEN_9657;
  wire [31:0] _GEN_9658;
  wire [31:0] _GEN_9659;
  wire [31:0] _GEN_9660;
  wire [31:0] _GEN_9661;
  wire [31:0] _GEN_9662;
  wire [31:0] _GEN_9663;
  wire [31:0] _GEN_9664;
  wire [31:0] _GEN_9665;
  wire [31:0] _GEN_9666;
  wire [31:0] _GEN_9667;
  wire [31:0] _GEN_9668;
  wire [31:0] _GEN_9669;
  wire [31:0] _GEN_9670;
  wire [31:0] _GEN_9671;
  wire [31:0] _GEN_9672;
  wire [31:0] _GEN_9673;
  wire [31:0] _GEN_9674;
  wire [31:0] _GEN_9675;
  wire [31:0] _GEN_9676;
  wire [31:0] _GEN_9677;
  wire [31:0] _GEN_9678;
  wire [31:0] _GEN_9679;
  wire [31:0] _GEN_9680;
  wire [31:0] _GEN_9681;
  wire [31:0] _GEN_9682;
  wire [31:0] _GEN_9683;
  wire [31:0] _GEN_9684;
  wire [31:0] _GEN_9685;
  wire [31:0] _GEN_9686;
  wire [31:0] _GEN_9687;
  wire [31:0] _GEN_9688;
  wire [31:0] _GEN_9689;
  wire [31:0] _GEN_9690;
  wire [31:0] _GEN_9691;
  wire [31:0] _GEN_9692;
  wire [31:0] _GEN_9693;
  wire [31:0] _GEN_9694;
  wire [31:0] _GEN_9695;
  wire [31:0] _GEN_9696;
  wire [31:0] _GEN_9697;
  wire [31:0] _GEN_9698;
  wire [31:0] _GEN_9699;
  wire [31:0] _GEN_9700;
  wire [31:0] _GEN_9701;
  wire [31:0] _GEN_9702;
  wire [31:0] _GEN_9703;
  wire [31:0] _GEN_9704;
  wire [31:0] _GEN_9705;
  wire [31:0] _GEN_9706;
  wire [31:0] _GEN_9707;
  wire [31:0] _GEN_9708;
  wire [31:0] _GEN_9709;
  wire [31:0] _GEN_9710;
  wire [31:0] _GEN_9711;
  wire [31:0] _GEN_9712;
  wire [31:0] _GEN_9713;
  wire [31:0] _GEN_9714;
  wire [31:0] _GEN_9715;
  wire [31:0] _GEN_9716;
  wire [31:0] _GEN_9717;
  wire [31:0] _GEN_9718;
  wire [31:0] _GEN_9719;
  wire [31:0] _GEN_9720;
  wire [31:0] _GEN_9721;
  wire [31:0] _GEN_9722;
  wire [31:0] _GEN_9723;
  wire [31:0] _GEN_9724;
  wire [31:0] _GEN_9725;
  wire [31:0] _GEN_9726;
  wire [31:0] _GEN_9727;
  wire [31:0] _GEN_9728;
  wire [31:0] _GEN_9729;
  wire [31:0] _GEN_9730;
  wire [31:0] _GEN_9731;
  wire [31:0] _GEN_9732;
  wire [31:0] _GEN_9733;
  wire [31:0] _GEN_9734;
  wire [31:0] _GEN_9735;
  wire [31:0] _GEN_9736;
  wire [31:0] _GEN_9737;
  wire [31:0] _GEN_9738;
  wire [31:0] _GEN_9739;
  wire [31:0] _GEN_9740;
  wire [31:0] _GEN_9741;
  wire [31:0] _GEN_9742;
  wire [31:0] _GEN_9743;
  wire [31:0] _GEN_9744;
  wire [31:0] _GEN_9745;
  wire [31:0] _GEN_9746;
  wire [31:0] _GEN_9747;
  wire [31:0] _GEN_9748;
  wire [31:0] _GEN_9749;
  wire [31:0] _GEN_9750;
  wire [31:0] _GEN_9751;
  wire [31:0] _GEN_9752;
  wire [31:0] _GEN_9753;
  wire [31:0] _GEN_9754;
  wire [31:0] _GEN_9755;
  wire [31:0] _GEN_9756;
  wire [31:0] _GEN_9757;
  wire [31:0] _GEN_9758;
  wire [31:0] _GEN_9759;
  wire [31:0] _GEN_9760;
  wire [31:0] _GEN_9761;
  wire [31:0] _GEN_9762;
  wire [31:0] _GEN_9763;
  wire [31:0] _GEN_9764;
  wire [31:0] _GEN_9765;
  wire [31:0] _GEN_9766;
  wire [31:0] _GEN_9767;
  wire [31:0] _GEN_9768;
  wire [31:0] _GEN_9769;
  wire [31:0] _GEN_9770;
  wire [31:0] _GEN_9771;
  wire [31:0] _GEN_9772;
  wire [31:0] _GEN_9773;
  wire [31:0] _GEN_9774;
  wire [31:0] _GEN_9775;
  wire [31:0] _GEN_9776;
  wire [31:0] _GEN_9777;
  wire [31:0] _GEN_9778;
  wire [31:0] _GEN_9779;
  wire [31:0] _GEN_9780;
  wire [31:0] _GEN_9781;
  wire [31:0] _GEN_9782;
  wire [31:0] _GEN_9783;
  wire [31:0] _GEN_9784;
  wire [31:0] _GEN_9785;
  wire [31:0] _GEN_9786;
  wire [31:0] _GEN_9787;
  wire [31:0] _GEN_9788;
  wire [31:0] _GEN_9789;
  wire [31:0] _GEN_9790;
  wire [31:0] _GEN_9791;
  wire [31:0] _GEN_9792;
  wire [31:0] _GEN_9793;
  wire [31:0] _GEN_9794;
  wire [31:0] _GEN_9795;
  wire [31:0] _GEN_9796;
  wire [31:0] _GEN_9797;
  wire [31:0] _GEN_9798;
  wire [31:0] _GEN_9799;
  wire [31:0] _GEN_9800;
  wire [31:0] _GEN_9801;
  wire [31:0] _GEN_9802;
  wire [31:0] _GEN_9803;
  wire [31:0] _GEN_9804;
  wire [31:0] _GEN_9805;
  wire [31:0] _GEN_9806;
  wire [31:0] _GEN_9807;
  wire [31:0] _GEN_9808;
  wire [31:0] _GEN_9809;
  wire [31:0] _GEN_9810;
  wire [31:0] _GEN_9811;
  wire [31:0] _GEN_9812;
  wire [31:0] _GEN_9813;
  wire [31:0] _GEN_9814;
  wire [31:0] _GEN_9815;
  wire [31:0] _GEN_9816;
  wire [31:0] _GEN_9817;
  wire [31:0] _GEN_9818;
  wire [31:0] _GEN_9819;
  wire [31:0] _GEN_9820;
  wire [31:0] _GEN_9821;
  wire [31:0] _GEN_9822;
  wire [31:0] _GEN_9823;
  wire [31:0] _GEN_9824;
  wire [31:0] _GEN_9825;
  wire [31:0] _GEN_9826;
  wire [31:0] _GEN_9827;
  wire [31:0] _GEN_9828;
  wire [31:0] _GEN_9829;
  wire [31:0] _GEN_9830;
  wire [31:0] _GEN_9831;
  wire [31:0] _GEN_9832;
  wire [31:0] _GEN_9833;
  wire [31:0] _GEN_9834;
  wire [31:0] _GEN_9835;
  wire [31:0] _GEN_9836;
  wire [31:0] _GEN_9837;
  wire [31:0] _GEN_9838;
  wire [31:0] _GEN_9839;
  wire [31:0] _GEN_9840;
  wire [31:0] _GEN_9841;
  wire [31:0] _GEN_9842;
  wire [31:0] _GEN_9843;
  wire [31:0] _GEN_9844;
  wire [31:0] _GEN_9845;
  wire [31:0] _GEN_9846;
  wire [31:0] _GEN_9847;
  wire [31:0] _GEN_9848;
  wire [31:0] _GEN_9849;
  wire [31:0] _GEN_9850;
  wire [31:0] _GEN_9851;
  wire [31:0] _GEN_9852;
  wire [31:0] _GEN_9853;
  wire [31:0] _GEN_9854;
  wire [31:0] _GEN_9855;
  wire [31:0] _GEN_9856;
  wire [31:0] _GEN_9857;
  wire [31:0] _GEN_9858;
  wire [31:0] _GEN_9859;
  wire [31:0] _GEN_9860;
  wire [31:0] _GEN_9861;
  wire [31:0] _GEN_9862;
  wire [31:0] _GEN_9863;
  wire [31:0] _GEN_9864;
  wire [31:0] _GEN_9865;
  wire [31:0] _GEN_9866;
  wire [31:0] _GEN_9867;
  wire [31:0] _GEN_9868;
  wire [31:0] _GEN_9869;
  wire [31:0] _GEN_9870;
  wire [31:0] _GEN_9871;
  wire [31:0] _GEN_9872;
  wire [31:0] _GEN_9873;
  wire [31:0] _GEN_9874;
  wire [31:0] _GEN_9875;
  wire [31:0] _GEN_9876;
  wire [31:0] _GEN_9877;
  wire [31:0] _GEN_9878;
  wire [31:0] _GEN_9879;
  wire [31:0] _GEN_9880;
  wire [31:0] _GEN_9881;
  wire [31:0] _GEN_9882;
  wire [31:0] _GEN_9883;
  wire [31:0] _GEN_9884;
  wire [31:0] _GEN_9885;
  wire [31:0] _GEN_9886;
  wire [31:0] _GEN_9887;
  wire [31:0] _GEN_9888;
  wire [31:0] _GEN_9889;
  wire [31:0] _GEN_9890;
  wire [31:0] _GEN_9891;
  wire [31:0] _GEN_9892;
  wire [31:0] _GEN_9893;
  wire [31:0] _GEN_9894;
  wire [31:0] _GEN_9895;
  wire [31:0] _GEN_9896;
  wire [31:0] _GEN_9897;
  wire [31:0] _GEN_9898;
  wire [31:0] _GEN_9899;
  wire [31:0] _GEN_9900;
  wire [31:0] _GEN_9901;
  wire [31:0] _GEN_9902;
  wire [31:0] _GEN_9903;
  wire [31:0] _GEN_9904;
  wire [31:0] _GEN_9905;
  wire [31:0] _GEN_9906;
  wire [31:0] _GEN_9907;
  wire [31:0] _GEN_9908;
  wire [31:0] _GEN_9909;
  wire [31:0] _GEN_9910;
  wire [31:0] _GEN_9911;
  wire [31:0] _GEN_9912;
  wire [31:0] _GEN_9913;
  wire [31:0] _GEN_9914;
  wire [31:0] _GEN_9915;
  wire [31:0] _GEN_9916;
  wire [31:0] _GEN_9917;
  wire [31:0] _GEN_9918;
  wire [31:0] _GEN_9919;
  wire [31:0] _GEN_9920;
  wire [31:0] _GEN_9921;
  wire [31:0] _GEN_9922;
  wire [31:0] _GEN_9923;
  wire [31:0] _GEN_9924;
  wire [31:0] _GEN_9925;
  wire [31:0] _GEN_9926;
  wire [31:0] _GEN_9927;
  wire [31:0] _GEN_9928;
  wire [31:0] _GEN_9929;
  wire [31:0] _GEN_9930;
  wire [31:0] _GEN_9931;
  wire [31:0] _GEN_9932;
  wire [31:0] _GEN_9933;
  wire [31:0] _GEN_9934;
  wire [31:0] _GEN_9935;
  wire [31:0] _GEN_9936;
  wire [31:0] _GEN_9937;
  wire [31:0] _GEN_9938;
  wire [31:0] _GEN_9939;
  wire [31:0] _GEN_9940;
  wire [31:0] _GEN_9941;
  wire [31:0] _GEN_9942;
  wire [31:0] _GEN_9943;
  wire [31:0] _GEN_9944;
  wire [31:0] _GEN_9945;
  wire [31:0] _GEN_9946;
  wire [31:0] _GEN_9947;
  wire [31:0] _GEN_9948;
  wire [31:0] _GEN_9949;
  wire [31:0] _GEN_9950;
  wire [31:0] _GEN_9951;
  wire [31:0] _GEN_9952;
  wire [31:0] _GEN_9953;
  wire [31:0] _GEN_9954;
  wire [31:0] _GEN_9955;
  wire [31:0] _GEN_9956;
  wire [31:0] _GEN_9957;
  wire [31:0] _GEN_9958;
  wire [31:0] _GEN_9959;
  wire [31:0] _GEN_9960;
  wire [31:0] _GEN_9961;
  wire [31:0] _GEN_9962;
  wire [31:0] _GEN_9963;
  wire [31:0] _GEN_9964;
  wire [31:0] _GEN_9965;
  wire [31:0] _GEN_9966;
  wire [31:0] _GEN_9967;
  wire [31:0] _GEN_9968;
  wire [31:0] _GEN_9969;
  wire [31:0] _GEN_9970;
  wire [31:0] _GEN_9971;
  wire [31:0] _GEN_9972;
  wire [31:0] _GEN_9973;
  wire [31:0] _GEN_9974;
  wire [31:0] _GEN_9975;
  wire [31:0] _GEN_9976;
  wire [31:0] _GEN_9977;
  wire [31:0] _GEN_9978;
  wire [31:0] _GEN_9979;
  wire [31:0] _GEN_9980;
  wire [31:0] _GEN_9981;
  wire [31:0] _GEN_9982;
  wire [31:0] _GEN_9983;
  wire [31:0] _GEN_9984;
  wire [31:0] _GEN_9985;
  wire [31:0] _GEN_9986;
  wire [31:0] _GEN_9987;
  wire [31:0] _GEN_9988;
  wire [31:0] _GEN_9989;
  wire [31:0] _GEN_9990;
  wire [31:0] _GEN_9991;
  wire [31:0] _GEN_9992;
  wire [31:0] _GEN_9993;
  wire [31:0] _GEN_9994;
  wire [31:0] _GEN_9995;
  wire [31:0] _GEN_9996;
  wire [31:0] _GEN_9997;
  wire [31:0] _GEN_9998;
  wire [31:0] _GEN_9999;
  wire [31:0] _GEN_10000;
  wire [31:0] _GEN_10001;
  wire [31:0] _GEN_10002;
  wire [31:0] _GEN_10003;
  wire [31:0] _GEN_10004;
  wire [31:0] _GEN_10005;
  wire [31:0] _GEN_10006;
  wire [31:0] _GEN_10007;
  wire [31:0] _GEN_10008;
  wire [31:0] _GEN_10009;
  wire [31:0] _GEN_10010;
  wire [31:0] _GEN_10011;
  wire [31:0] _GEN_10012;
  wire [31:0] _GEN_10013;
  wire [31:0] _GEN_10014;
  wire [31:0] _GEN_10015;
  wire [31:0] _GEN_10016;
  wire [31:0] _GEN_10017;
  wire [31:0] _GEN_10018;
  wire [31:0] _GEN_10019;
  wire [31:0] _GEN_10020;
  wire [31:0] _GEN_10021;
  wire [31:0] _GEN_10022;
  wire [31:0] _GEN_10023;
  wire [31:0] _GEN_10024;
  wire [31:0] _GEN_10025;
  wire [31:0] _GEN_10026;
  wire [31:0] _GEN_10027;
  wire [31:0] _GEN_10028;
  wire [31:0] _GEN_10029;
  wire [31:0] _GEN_10030;
  wire [31:0] _GEN_10031;
  wire [31:0] _GEN_10032;
  wire [31:0] _GEN_10033;
  wire [31:0] _GEN_10034;
  wire [31:0] _GEN_10035;
  wire [31:0] _GEN_10036;
  wire [31:0] _GEN_10037;
  wire [31:0] _GEN_10038;
  wire [31:0] _GEN_10039;
  wire [31:0] _GEN_10040;
  wire [31:0] _GEN_10041;
  wire [31:0] _GEN_10042;
  wire [31:0] _GEN_10043;
  wire [31:0] _GEN_10044;
  wire [31:0] _GEN_10045;
  wire [31:0] _GEN_10046;
  wire [31:0] _GEN_10047;
  wire [31:0] _GEN_10048;
  wire [31:0] _GEN_10049;
  wire [31:0] _GEN_10050;
  wire [31:0] _GEN_10051;
  wire [31:0] _GEN_10052;
  wire [31:0] _GEN_10053;
  wire [31:0] _GEN_10054;
  wire [31:0] _GEN_10055;
  wire [31:0] _GEN_10056;
  wire [31:0] _GEN_10057;
  wire [31:0] _GEN_10058;
  wire [31:0] _GEN_10059;
  wire [31:0] _GEN_10060;
  wire [31:0] _GEN_10061;
  wire [31:0] _GEN_10062;
  wire [31:0] _GEN_10063;
  wire [31:0] _GEN_10064;
  wire [31:0] _GEN_10065;
  wire [31:0] _GEN_10066;
  wire [31:0] _GEN_10067;
  wire [31:0] _GEN_10068;
  wire [31:0] _GEN_10069;
  wire [31:0] _GEN_10070;
  wire [31:0] _GEN_10071;
  wire [31:0] _GEN_10072;
  wire [31:0] _GEN_10073;
  wire [31:0] _GEN_10074;
  wire [31:0] _GEN_10075;
  wire [31:0] _GEN_10076;
  wire [31:0] _GEN_10077;
  wire [31:0] _GEN_10078;
  wire [31:0] _GEN_10079;
  wire [31:0] _GEN_10080;
  wire [31:0] _GEN_10081;
  wire [31:0] _GEN_10082;
  wire [31:0] _GEN_10083;
  wire [31:0] _GEN_10084;
  wire [31:0] _GEN_10085;
  wire [31:0] _GEN_10086;
  wire [31:0] _GEN_10087;
  wire [31:0] _GEN_10088;
  wire [31:0] _GEN_10089;
  wire [31:0] _GEN_10090;
  wire [31:0] _GEN_10091;
  wire [31:0] _GEN_10092;
  wire [31:0] _GEN_10093;
  wire [31:0] _GEN_10094;
  wire [31:0] _GEN_10095;
  wire [31:0] _GEN_10096;
  wire [31:0] _GEN_10097;
  wire [31:0] _GEN_10098;
  wire [31:0] _GEN_10099;
  wire [31:0] _GEN_10100;
  wire [31:0] _GEN_10101;
  wire [31:0] _GEN_10102;
  wire [31:0] _GEN_10103;
  wire [31:0] _GEN_10104;
  wire [31:0] _GEN_10105;
  wire [31:0] _GEN_10106;
  wire [31:0] _GEN_10107;
  wire [31:0] _GEN_10108;
  wire [31:0] _GEN_10109;
  wire [31:0] _GEN_10110;
  wire [31:0] _GEN_10111;
  wire [31:0] _GEN_10112;
  wire [31:0] _GEN_10113;
  wire [31:0] _GEN_10114;
  wire [31:0] _GEN_10115;
  wire [31:0] _GEN_10116;
  wire [31:0] _GEN_10117;
  wire [31:0] _GEN_10118;
  wire [31:0] _GEN_10119;
  wire [31:0] _GEN_10120;
  wire [31:0] _GEN_10121;
  wire [31:0] _GEN_10122;
  wire [31:0] _GEN_10123;
  wire [31:0] _GEN_10124;
  wire [31:0] _GEN_10125;
  wire [31:0] _GEN_10126;
  wire [31:0] _GEN_10127;
  wire [31:0] _GEN_10128;
  wire [31:0] _GEN_10129;
  wire [31:0] _GEN_10130;
  wire [31:0] _GEN_10131;
  wire [31:0] _GEN_10132;
  wire [31:0] _GEN_10133;
  wire [31:0] _GEN_10134;
  wire [31:0] _GEN_10135;
  wire [31:0] _GEN_10136;
  wire [31:0] _GEN_10137;
  wire [31:0] _GEN_10138;
  wire [31:0] _GEN_10139;
  wire [31:0] _GEN_10140;
  wire [31:0] _GEN_10141;
  wire [31:0] _GEN_10142;
  wire [31:0] _GEN_10143;
  wire [31:0] _GEN_10144;
  wire [31:0] _GEN_10145;
  wire [31:0] _GEN_10146;
  wire [31:0] _GEN_10147;
  wire [31:0] _GEN_10148;
  wire [31:0] _GEN_10149;
  wire [31:0] _GEN_10150;
  wire [31:0] _GEN_10151;
  wire [31:0] _GEN_10152;
  wire [31:0] _GEN_10153;
  wire [31:0] _GEN_10154;
  wire [31:0] _GEN_10155;
  wire [31:0] _GEN_10156;
  wire [31:0] _GEN_10157;
  wire [31:0] _GEN_10158;
  wire [31:0] _GEN_10159;
  wire [31:0] _GEN_10160;
  wire [31:0] _GEN_10161;
  wire [31:0] _GEN_10162;
  wire [31:0] _GEN_10163;
  wire [31:0] _GEN_10164;
  wire [31:0] _GEN_10165;
  wire [31:0] _GEN_10166;
  wire [31:0] _GEN_10167;
  wire [31:0] _GEN_10168;
  wire [31:0] _GEN_10169;
  wire [31:0] _GEN_10170;
  wire [31:0] _GEN_10171;
  wire [31:0] _GEN_10172;
  wire [31:0] _GEN_10173;
  wire [31:0] _GEN_10174;
  wire [31:0] _GEN_10175;
  wire [31:0] _GEN_10176;
  wire [31:0] _GEN_10177;
  wire [31:0] _GEN_10178;
  wire [31:0] _GEN_10179;
  wire [31:0] _GEN_10180;
  wire [31:0] _GEN_10181;
  wire [31:0] _GEN_10182;
  wire [31:0] _GEN_10183;
  wire [31:0] _GEN_10184;
  wire [31:0] _GEN_10185;
  wire [31:0] _GEN_10186;
  wire [31:0] _GEN_10187;
  wire [31:0] _GEN_10188;
  wire [31:0] _GEN_10189;
  wire [31:0] _GEN_10190;
  wire [31:0] _GEN_10191;
  wire [31:0] _GEN_10192;
  wire [31:0] _GEN_10193;
  wire [31:0] _GEN_10194;
  wire [31:0] _GEN_10195;
  wire [31:0] _GEN_10196;
  wire [31:0] _GEN_10197;
  wire [31:0] _GEN_10198;
  wire [31:0] _GEN_10199;
  wire [31:0] _GEN_10200;
  wire [31:0] _GEN_10201;
  wire [31:0] _GEN_10202;
  wire [31:0] _GEN_10203;
  wire [31:0] _GEN_10204;
  wire [31:0] _GEN_10205;
  wire [31:0] _GEN_10206;
  wire [31:0] _GEN_10207;
  wire [31:0] _GEN_10208;
  wire [31:0] _GEN_10209;
  wire [31:0] _GEN_10210;
  wire [31:0] _GEN_10211;
  wire [31:0] _GEN_10212;
  wire [31:0] _GEN_10213;
  wire [31:0] _GEN_10214;
  wire [31:0] _GEN_10215;
  wire [31:0] _GEN_10216;
  wire [31:0] _GEN_10217;
  wire [31:0] _GEN_10218;
  wire [31:0] _GEN_10219;
  wire [31:0] _GEN_10220;
  wire [31:0] _GEN_10221;
  wire [31:0] _GEN_10222;
  wire [31:0] _GEN_10223;
  wire [31:0] _GEN_10224;
  wire [31:0] _GEN_10225;
  wire [31:0] _GEN_10226;
  wire [31:0] _GEN_10227;
  wire [31:0] _GEN_10228;
  wire [31:0] _GEN_10229;
  wire [31:0] _GEN_10230;
  wire [31:0] _GEN_10231;
  wire [31:0] _GEN_10232;
  wire [31:0] _GEN_10233;
  wire [31:0] _GEN_10234;
  wire [31:0] _GEN_10235;
  wire [31:0] _GEN_10236;
  wire [31:0] _GEN_10237;
  wire [31:0] _GEN_10238;
  wire [31:0] _GEN_10239;
  wire [31:0] _GEN_10240;
  wire [31:0] _GEN_10241;
  wire [31:0] _GEN_10242;
  wire [31:0] _GEN_10243;
  wire [31:0] _GEN_10244;
  wire [31:0] _GEN_10245;
  wire [31:0] _GEN_5;
  assign _T_12316 = wen[0];
  assign _T_12319 = wdata[7:0];
  assign _T_12323 = addr[10:0];
  assign _GEN_6 = 11'h1 == _T_12323 ? mem_1 : mem_0;
  assign _GEN_7 = 11'h2 == _T_12323 ? mem_2 : _GEN_6;
  assign _GEN_8 = 11'h3 == _T_12323 ? mem_3 : _GEN_7;
  assign _GEN_9 = 11'h4 == _T_12323 ? mem_4 : _GEN_8;
  assign _GEN_10 = 11'h5 == _T_12323 ? mem_5 : _GEN_9;
  assign _GEN_11 = 11'h6 == _T_12323 ? mem_6 : _GEN_10;
  assign _GEN_12 = 11'h7 == _T_12323 ? mem_7 : _GEN_11;
  assign _GEN_13 = 11'h8 == _T_12323 ? mem_8 : _GEN_12;
  assign _GEN_14 = 11'h9 == _T_12323 ? mem_9 : _GEN_13;
  assign _GEN_15 = 11'ha == _T_12323 ? mem_10 : _GEN_14;
  assign _GEN_16 = 11'hb == _T_12323 ? mem_11 : _GEN_15;
  assign _GEN_17 = 11'hc == _T_12323 ? mem_12 : _GEN_16;
  assign _GEN_18 = 11'hd == _T_12323 ? mem_13 : _GEN_17;
  assign _GEN_19 = 11'he == _T_12323 ? mem_14 : _GEN_18;
  assign _GEN_20 = 11'hf == _T_12323 ? mem_15 : _GEN_19;
  assign _GEN_21 = 11'h10 == _T_12323 ? mem_16 : _GEN_20;
  assign _GEN_22 = 11'h11 == _T_12323 ? mem_17 : _GEN_21;
  assign _GEN_23 = 11'h12 == _T_12323 ? mem_18 : _GEN_22;
  assign _GEN_24 = 11'h13 == _T_12323 ? mem_19 : _GEN_23;
  assign _GEN_25 = 11'h14 == _T_12323 ? mem_20 : _GEN_24;
  assign _GEN_26 = 11'h15 == _T_12323 ? mem_21 : _GEN_25;
  assign _GEN_27 = 11'h16 == _T_12323 ? mem_22 : _GEN_26;
  assign _GEN_28 = 11'h17 == _T_12323 ? mem_23 : _GEN_27;
  assign _GEN_29 = 11'h18 == _T_12323 ? mem_24 : _GEN_28;
  assign _GEN_30 = 11'h19 == _T_12323 ? mem_25 : _GEN_29;
  assign _GEN_31 = 11'h1a == _T_12323 ? mem_26 : _GEN_30;
  assign _GEN_32 = 11'h1b == _T_12323 ? mem_27 : _GEN_31;
  assign _GEN_33 = 11'h1c == _T_12323 ? mem_28 : _GEN_32;
  assign _GEN_34 = 11'h1d == _T_12323 ? mem_29 : _GEN_33;
  assign _GEN_35 = 11'h1e == _T_12323 ? mem_30 : _GEN_34;
  assign _GEN_36 = 11'h1f == _T_12323 ? mem_31 : _GEN_35;
  assign _GEN_37 = 11'h20 == _T_12323 ? mem_32 : _GEN_36;
  assign _GEN_38 = 11'h21 == _T_12323 ? mem_33 : _GEN_37;
  assign _GEN_39 = 11'h22 == _T_12323 ? mem_34 : _GEN_38;
  assign _GEN_40 = 11'h23 == _T_12323 ? mem_35 : _GEN_39;
  assign _GEN_41 = 11'h24 == _T_12323 ? mem_36 : _GEN_40;
  assign _GEN_42 = 11'h25 == _T_12323 ? mem_37 : _GEN_41;
  assign _GEN_43 = 11'h26 == _T_12323 ? mem_38 : _GEN_42;
  assign _GEN_44 = 11'h27 == _T_12323 ? mem_39 : _GEN_43;
  assign _GEN_45 = 11'h28 == _T_12323 ? mem_40 : _GEN_44;
  assign _GEN_46 = 11'h29 == _T_12323 ? mem_41 : _GEN_45;
  assign _GEN_47 = 11'h2a == _T_12323 ? mem_42 : _GEN_46;
  assign _GEN_48 = 11'h2b == _T_12323 ? mem_43 : _GEN_47;
  assign _GEN_49 = 11'h2c == _T_12323 ? mem_44 : _GEN_48;
  assign _GEN_50 = 11'h2d == _T_12323 ? mem_45 : _GEN_49;
  assign _GEN_51 = 11'h2e == _T_12323 ? mem_46 : _GEN_50;
  assign _GEN_52 = 11'h2f == _T_12323 ? mem_47 : _GEN_51;
  assign _GEN_53 = 11'h30 == _T_12323 ? mem_48 : _GEN_52;
  assign _GEN_54 = 11'h31 == _T_12323 ? mem_49 : _GEN_53;
  assign _GEN_55 = 11'h32 == _T_12323 ? mem_50 : _GEN_54;
  assign _GEN_56 = 11'h33 == _T_12323 ? mem_51 : _GEN_55;
  assign _GEN_57 = 11'h34 == _T_12323 ? mem_52 : _GEN_56;
  assign _GEN_58 = 11'h35 == _T_12323 ? mem_53 : _GEN_57;
  assign _GEN_59 = 11'h36 == _T_12323 ? mem_54 : _GEN_58;
  assign _GEN_60 = 11'h37 == _T_12323 ? mem_55 : _GEN_59;
  assign _GEN_61 = 11'h38 == _T_12323 ? mem_56 : _GEN_60;
  assign _GEN_62 = 11'h39 == _T_12323 ? mem_57 : _GEN_61;
  assign _GEN_63 = 11'h3a == _T_12323 ? mem_58 : _GEN_62;
  assign _GEN_64 = 11'h3b == _T_12323 ? mem_59 : _GEN_63;
  assign _GEN_65 = 11'h3c == _T_12323 ? mem_60 : _GEN_64;
  assign _GEN_66 = 11'h3d == _T_12323 ? mem_61 : _GEN_65;
  assign _GEN_67 = 11'h3e == _T_12323 ? mem_62 : _GEN_66;
  assign _GEN_68 = 11'h3f == _T_12323 ? mem_63 : _GEN_67;
  assign _GEN_69 = 11'h40 == _T_12323 ? mem_64 : _GEN_68;
  assign _GEN_70 = 11'h41 == _T_12323 ? mem_65 : _GEN_69;
  assign _GEN_71 = 11'h42 == _T_12323 ? mem_66 : _GEN_70;
  assign _GEN_72 = 11'h43 == _T_12323 ? mem_67 : _GEN_71;
  assign _GEN_73 = 11'h44 == _T_12323 ? mem_68 : _GEN_72;
  assign _GEN_74 = 11'h45 == _T_12323 ? mem_69 : _GEN_73;
  assign _GEN_75 = 11'h46 == _T_12323 ? mem_70 : _GEN_74;
  assign _GEN_76 = 11'h47 == _T_12323 ? mem_71 : _GEN_75;
  assign _GEN_77 = 11'h48 == _T_12323 ? mem_72 : _GEN_76;
  assign _GEN_78 = 11'h49 == _T_12323 ? mem_73 : _GEN_77;
  assign _GEN_79 = 11'h4a == _T_12323 ? mem_74 : _GEN_78;
  assign _GEN_80 = 11'h4b == _T_12323 ? mem_75 : _GEN_79;
  assign _GEN_81 = 11'h4c == _T_12323 ? mem_76 : _GEN_80;
  assign _GEN_82 = 11'h4d == _T_12323 ? mem_77 : _GEN_81;
  assign _GEN_83 = 11'h4e == _T_12323 ? mem_78 : _GEN_82;
  assign _GEN_84 = 11'h4f == _T_12323 ? mem_79 : _GEN_83;
  assign _GEN_85 = 11'h50 == _T_12323 ? mem_80 : _GEN_84;
  assign _GEN_86 = 11'h51 == _T_12323 ? mem_81 : _GEN_85;
  assign _GEN_87 = 11'h52 == _T_12323 ? mem_82 : _GEN_86;
  assign _GEN_88 = 11'h53 == _T_12323 ? mem_83 : _GEN_87;
  assign _GEN_89 = 11'h54 == _T_12323 ? mem_84 : _GEN_88;
  assign _GEN_90 = 11'h55 == _T_12323 ? mem_85 : _GEN_89;
  assign _GEN_91 = 11'h56 == _T_12323 ? mem_86 : _GEN_90;
  assign _GEN_92 = 11'h57 == _T_12323 ? mem_87 : _GEN_91;
  assign _GEN_93 = 11'h58 == _T_12323 ? mem_88 : _GEN_92;
  assign _GEN_94 = 11'h59 == _T_12323 ? mem_89 : _GEN_93;
  assign _GEN_95 = 11'h5a == _T_12323 ? mem_90 : _GEN_94;
  assign _GEN_96 = 11'h5b == _T_12323 ? mem_91 : _GEN_95;
  assign _GEN_97 = 11'h5c == _T_12323 ? mem_92 : _GEN_96;
  assign _GEN_98 = 11'h5d == _T_12323 ? mem_93 : _GEN_97;
  assign _GEN_99 = 11'h5e == _T_12323 ? mem_94 : _GEN_98;
  assign _GEN_100 = 11'h5f == _T_12323 ? mem_95 : _GEN_99;
  assign _GEN_101 = 11'h60 == _T_12323 ? mem_96 : _GEN_100;
  assign _GEN_102 = 11'h61 == _T_12323 ? mem_97 : _GEN_101;
  assign _GEN_103 = 11'h62 == _T_12323 ? mem_98 : _GEN_102;
  assign _GEN_104 = 11'h63 == _T_12323 ? mem_99 : _GEN_103;
  assign _GEN_105 = 11'h64 == _T_12323 ? mem_100 : _GEN_104;
  assign _GEN_106 = 11'h65 == _T_12323 ? mem_101 : _GEN_105;
  assign _GEN_107 = 11'h66 == _T_12323 ? mem_102 : _GEN_106;
  assign _GEN_108 = 11'h67 == _T_12323 ? mem_103 : _GEN_107;
  assign _GEN_109 = 11'h68 == _T_12323 ? mem_104 : _GEN_108;
  assign _GEN_110 = 11'h69 == _T_12323 ? mem_105 : _GEN_109;
  assign _GEN_111 = 11'h6a == _T_12323 ? mem_106 : _GEN_110;
  assign _GEN_112 = 11'h6b == _T_12323 ? mem_107 : _GEN_111;
  assign _GEN_113 = 11'h6c == _T_12323 ? mem_108 : _GEN_112;
  assign _GEN_114 = 11'h6d == _T_12323 ? mem_109 : _GEN_113;
  assign _GEN_115 = 11'h6e == _T_12323 ? mem_110 : _GEN_114;
  assign _GEN_116 = 11'h6f == _T_12323 ? mem_111 : _GEN_115;
  assign _GEN_117 = 11'h70 == _T_12323 ? mem_112 : _GEN_116;
  assign _GEN_118 = 11'h71 == _T_12323 ? mem_113 : _GEN_117;
  assign _GEN_119 = 11'h72 == _T_12323 ? mem_114 : _GEN_118;
  assign _GEN_120 = 11'h73 == _T_12323 ? mem_115 : _GEN_119;
  assign _GEN_121 = 11'h74 == _T_12323 ? mem_116 : _GEN_120;
  assign _GEN_122 = 11'h75 == _T_12323 ? mem_117 : _GEN_121;
  assign _GEN_123 = 11'h76 == _T_12323 ? mem_118 : _GEN_122;
  assign _GEN_124 = 11'h77 == _T_12323 ? mem_119 : _GEN_123;
  assign _GEN_125 = 11'h78 == _T_12323 ? mem_120 : _GEN_124;
  assign _GEN_126 = 11'h79 == _T_12323 ? mem_121 : _GEN_125;
  assign _GEN_127 = 11'h7a == _T_12323 ? mem_122 : _GEN_126;
  assign _GEN_128 = 11'h7b == _T_12323 ? mem_123 : _GEN_127;
  assign _GEN_129 = 11'h7c == _T_12323 ? mem_124 : _GEN_128;
  assign _GEN_130 = 11'h7d == _T_12323 ? mem_125 : _GEN_129;
  assign _GEN_131 = 11'h7e == _T_12323 ? mem_126 : _GEN_130;
  assign _GEN_132 = 11'h7f == _T_12323 ? mem_127 : _GEN_131;
  assign _GEN_133 = 11'h80 == _T_12323 ? mem_128 : _GEN_132;
  assign _GEN_134 = 11'h81 == _T_12323 ? mem_129 : _GEN_133;
  assign _GEN_135 = 11'h82 == _T_12323 ? mem_130 : _GEN_134;
  assign _GEN_136 = 11'h83 == _T_12323 ? mem_131 : _GEN_135;
  assign _GEN_137 = 11'h84 == _T_12323 ? mem_132 : _GEN_136;
  assign _GEN_138 = 11'h85 == _T_12323 ? mem_133 : _GEN_137;
  assign _GEN_139 = 11'h86 == _T_12323 ? mem_134 : _GEN_138;
  assign _GEN_140 = 11'h87 == _T_12323 ? mem_135 : _GEN_139;
  assign _GEN_141 = 11'h88 == _T_12323 ? mem_136 : _GEN_140;
  assign _GEN_142 = 11'h89 == _T_12323 ? mem_137 : _GEN_141;
  assign _GEN_143 = 11'h8a == _T_12323 ? mem_138 : _GEN_142;
  assign _GEN_144 = 11'h8b == _T_12323 ? mem_139 : _GEN_143;
  assign _GEN_145 = 11'h8c == _T_12323 ? mem_140 : _GEN_144;
  assign _GEN_146 = 11'h8d == _T_12323 ? mem_141 : _GEN_145;
  assign _GEN_147 = 11'h8e == _T_12323 ? mem_142 : _GEN_146;
  assign _GEN_148 = 11'h8f == _T_12323 ? mem_143 : _GEN_147;
  assign _GEN_149 = 11'h90 == _T_12323 ? mem_144 : _GEN_148;
  assign _GEN_150 = 11'h91 == _T_12323 ? mem_145 : _GEN_149;
  assign _GEN_151 = 11'h92 == _T_12323 ? mem_146 : _GEN_150;
  assign _GEN_152 = 11'h93 == _T_12323 ? mem_147 : _GEN_151;
  assign _GEN_153 = 11'h94 == _T_12323 ? mem_148 : _GEN_152;
  assign _GEN_154 = 11'h95 == _T_12323 ? mem_149 : _GEN_153;
  assign _GEN_155 = 11'h96 == _T_12323 ? mem_150 : _GEN_154;
  assign _GEN_156 = 11'h97 == _T_12323 ? mem_151 : _GEN_155;
  assign _GEN_157 = 11'h98 == _T_12323 ? mem_152 : _GEN_156;
  assign _GEN_158 = 11'h99 == _T_12323 ? mem_153 : _GEN_157;
  assign _GEN_159 = 11'h9a == _T_12323 ? mem_154 : _GEN_158;
  assign _GEN_160 = 11'h9b == _T_12323 ? mem_155 : _GEN_159;
  assign _GEN_161 = 11'h9c == _T_12323 ? mem_156 : _GEN_160;
  assign _GEN_162 = 11'h9d == _T_12323 ? mem_157 : _GEN_161;
  assign _GEN_163 = 11'h9e == _T_12323 ? mem_158 : _GEN_162;
  assign _GEN_164 = 11'h9f == _T_12323 ? mem_159 : _GEN_163;
  assign _GEN_165 = 11'ha0 == _T_12323 ? mem_160 : _GEN_164;
  assign _GEN_166 = 11'ha1 == _T_12323 ? mem_161 : _GEN_165;
  assign _GEN_167 = 11'ha2 == _T_12323 ? mem_162 : _GEN_166;
  assign _GEN_168 = 11'ha3 == _T_12323 ? mem_163 : _GEN_167;
  assign _GEN_169 = 11'ha4 == _T_12323 ? mem_164 : _GEN_168;
  assign _GEN_170 = 11'ha5 == _T_12323 ? mem_165 : _GEN_169;
  assign _GEN_171 = 11'ha6 == _T_12323 ? mem_166 : _GEN_170;
  assign _GEN_172 = 11'ha7 == _T_12323 ? mem_167 : _GEN_171;
  assign _GEN_173 = 11'ha8 == _T_12323 ? mem_168 : _GEN_172;
  assign _GEN_174 = 11'ha9 == _T_12323 ? mem_169 : _GEN_173;
  assign _GEN_175 = 11'haa == _T_12323 ? mem_170 : _GEN_174;
  assign _GEN_176 = 11'hab == _T_12323 ? mem_171 : _GEN_175;
  assign _GEN_177 = 11'hac == _T_12323 ? mem_172 : _GEN_176;
  assign _GEN_178 = 11'had == _T_12323 ? mem_173 : _GEN_177;
  assign _GEN_179 = 11'hae == _T_12323 ? mem_174 : _GEN_178;
  assign _GEN_180 = 11'haf == _T_12323 ? mem_175 : _GEN_179;
  assign _GEN_181 = 11'hb0 == _T_12323 ? mem_176 : _GEN_180;
  assign _GEN_182 = 11'hb1 == _T_12323 ? mem_177 : _GEN_181;
  assign _GEN_183 = 11'hb2 == _T_12323 ? mem_178 : _GEN_182;
  assign _GEN_184 = 11'hb3 == _T_12323 ? mem_179 : _GEN_183;
  assign _GEN_185 = 11'hb4 == _T_12323 ? mem_180 : _GEN_184;
  assign _GEN_186 = 11'hb5 == _T_12323 ? mem_181 : _GEN_185;
  assign _GEN_187 = 11'hb6 == _T_12323 ? mem_182 : _GEN_186;
  assign _GEN_188 = 11'hb7 == _T_12323 ? mem_183 : _GEN_187;
  assign _GEN_189 = 11'hb8 == _T_12323 ? mem_184 : _GEN_188;
  assign _GEN_190 = 11'hb9 == _T_12323 ? mem_185 : _GEN_189;
  assign _GEN_191 = 11'hba == _T_12323 ? mem_186 : _GEN_190;
  assign _GEN_192 = 11'hbb == _T_12323 ? mem_187 : _GEN_191;
  assign _GEN_193 = 11'hbc == _T_12323 ? mem_188 : _GEN_192;
  assign _GEN_194 = 11'hbd == _T_12323 ? mem_189 : _GEN_193;
  assign _GEN_195 = 11'hbe == _T_12323 ? mem_190 : _GEN_194;
  assign _GEN_196 = 11'hbf == _T_12323 ? mem_191 : _GEN_195;
  assign _GEN_197 = 11'hc0 == _T_12323 ? mem_192 : _GEN_196;
  assign _GEN_198 = 11'hc1 == _T_12323 ? mem_193 : _GEN_197;
  assign _GEN_199 = 11'hc2 == _T_12323 ? mem_194 : _GEN_198;
  assign _GEN_200 = 11'hc3 == _T_12323 ? mem_195 : _GEN_199;
  assign _GEN_201 = 11'hc4 == _T_12323 ? mem_196 : _GEN_200;
  assign _GEN_202 = 11'hc5 == _T_12323 ? mem_197 : _GEN_201;
  assign _GEN_203 = 11'hc6 == _T_12323 ? mem_198 : _GEN_202;
  assign _GEN_204 = 11'hc7 == _T_12323 ? mem_199 : _GEN_203;
  assign _GEN_205 = 11'hc8 == _T_12323 ? mem_200 : _GEN_204;
  assign _GEN_206 = 11'hc9 == _T_12323 ? mem_201 : _GEN_205;
  assign _GEN_207 = 11'hca == _T_12323 ? mem_202 : _GEN_206;
  assign _GEN_208 = 11'hcb == _T_12323 ? mem_203 : _GEN_207;
  assign _GEN_209 = 11'hcc == _T_12323 ? mem_204 : _GEN_208;
  assign _GEN_210 = 11'hcd == _T_12323 ? mem_205 : _GEN_209;
  assign _GEN_211 = 11'hce == _T_12323 ? mem_206 : _GEN_210;
  assign _GEN_212 = 11'hcf == _T_12323 ? mem_207 : _GEN_211;
  assign _GEN_213 = 11'hd0 == _T_12323 ? mem_208 : _GEN_212;
  assign _GEN_214 = 11'hd1 == _T_12323 ? mem_209 : _GEN_213;
  assign _GEN_215 = 11'hd2 == _T_12323 ? mem_210 : _GEN_214;
  assign _GEN_216 = 11'hd3 == _T_12323 ? mem_211 : _GEN_215;
  assign _GEN_217 = 11'hd4 == _T_12323 ? mem_212 : _GEN_216;
  assign _GEN_218 = 11'hd5 == _T_12323 ? mem_213 : _GEN_217;
  assign _GEN_219 = 11'hd6 == _T_12323 ? mem_214 : _GEN_218;
  assign _GEN_220 = 11'hd7 == _T_12323 ? mem_215 : _GEN_219;
  assign _GEN_221 = 11'hd8 == _T_12323 ? mem_216 : _GEN_220;
  assign _GEN_222 = 11'hd9 == _T_12323 ? mem_217 : _GEN_221;
  assign _GEN_223 = 11'hda == _T_12323 ? mem_218 : _GEN_222;
  assign _GEN_224 = 11'hdb == _T_12323 ? mem_219 : _GEN_223;
  assign _GEN_225 = 11'hdc == _T_12323 ? mem_220 : _GEN_224;
  assign _GEN_226 = 11'hdd == _T_12323 ? mem_221 : _GEN_225;
  assign _GEN_227 = 11'hde == _T_12323 ? mem_222 : _GEN_226;
  assign _GEN_228 = 11'hdf == _T_12323 ? mem_223 : _GEN_227;
  assign _GEN_229 = 11'he0 == _T_12323 ? mem_224 : _GEN_228;
  assign _GEN_230 = 11'he1 == _T_12323 ? mem_225 : _GEN_229;
  assign _GEN_231 = 11'he2 == _T_12323 ? mem_226 : _GEN_230;
  assign _GEN_232 = 11'he3 == _T_12323 ? mem_227 : _GEN_231;
  assign _GEN_233 = 11'he4 == _T_12323 ? mem_228 : _GEN_232;
  assign _GEN_234 = 11'he5 == _T_12323 ? mem_229 : _GEN_233;
  assign _GEN_235 = 11'he6 == _T_12323 ? mem_230 : _GEN_234;
  assign _GEN_236 = 11'he7 == _T_12323 ? mem_231 : _GEN_235;
  assign _GEN_237 = 11'he8 == _T_12323 ? mem_232 : _GEN_236;
  assign _GEN_238 = 11'he9 == _T_12323 ? mem_233 : _GEN_237;
  assign _GEN_239 = 11'hea == _T_12323 ? mem_234 : _GEN_238;
  assign _GEN_240 = 11'heb == _T_12323 ? mem_235 : _GEN_239;
  assign _GEN_241 = 11'hec == _T_12323 ? mem_236 : _GEN_240;
  assign _GEN_242 = 11'hed == _T_12323 ? mem_237 : _GEN_241;
  assign _GEN_243 = 11'hee == _T_12323 ? mem_238 : _GEN_242;
  assign _GEN_244 = 11'hef == _T_12323 ? mem_239 : _GEN_243;
  assign _GEN_245 = 11'hf0 == _T_12323 ? mem_240 : _GEN_244;
  assign _GEN_246 = 11'hf1 == _T_12323 ? mem_241 : _GEN_245;
  assign _GEN_247 = 11'hf2 == _T_12323 ? mem_242 : _GEN_246;
  assign _GEN_248 = 11'hf3 == _T_12323 ? mem_243 : _GEN_247;
  assign _GEN_249 = 11'hf4 == _T_12323 ? mem_244 : _GEN_248;
  assign _GEN_250 = 11'hf5 == _T_12323 ? mem_245 : _GEN_249;
  assign _GEN_251 = 11'hf6 == _T_12323 ? mem_246 : _GEN_250;
  assign _GEN_252 = 11'hf7 == _T_12323 ? mem_247 : _GEN_251;
  assign _GEN_253 = 11'hf8 == _T_12323 ? mem_248 : _GEN_252;
  assign _GEN_254 = 11'hf9 == _T_12323 ? mem_249 : _GEN_253;
  assign _GEN_255 = 11'hfa == _T_12323 ? mem_250 : _GEN_254;
  assign _GEN_256 = 11'hfb == _T_12323 ? mem_251 : _GEN_255;
  assign _GEN_257 = 11'hfc == _T_12323 ? mem_252 : _GEN_256;
  assign _GEN_258 = 11'hfd == _T_12323 ? mem_253 : _GEN_257;
  assign _GEN_259 = 11'hfe == _T_12323 ? mem_254 : _GEN_258;
  assign _GEN_260 = 11'hff == _T_12323 ? mem_255 : _GEN_259;
  assign _GEN_261 = 11'h100 == _T_12323 ? mem_256 : _GEN_260;
  assign _GEN_262 = 11'h101 == _T_12323 ? mem_257 : _GEN_261;
  assign _GEN_263 = 11'h102 == _T_12323 ? mem_258 : _GEN_262;
  assign _GEN_264 = 11'h103 == _T_12323 ? mem_259 : _GEN_263;
  assign _GEN_265 = 11'h104 == _T_12323 ? mem_260 : _GEN_264;
  assign _GEN_266 = 11'h105 == _T_12323 ? mem_261 : _GEN_265;
  assign _GEN_267 = 11'h106 == _T_12323 ? mem_262 : _GEN_266;
  assign _GEN_268 = 11'h107 == _T_12323 ? mem_263 : _GEN_267;
  assign _GEN_269 = 11'h108 == _T_12323 ? mem_264 : _GEN_268;
  assign _GEN_270 = 11'h109 == _T_12323 ? mem_265 : _GEN_269;
  assign _GEN_271 = 11'h10a == _T_12323 ? mem_266 : _GEN_270;
  assign _GEN_272 = 11'h10b == _T_12323 ? mem_267 : _GEN_271;
  assign _GEN_273 = 11'h10c == _T_12323 ? mem_268 : _GEN_272;
  assign _GEN_274 = 11'h10d == _T_12323 ? mem_269 : _GEN_273;
  assign _GEN_275 = 11'h10e == _T_12323 ? mem_270 : _GEN_274;
  assign _GEN_276 = 11'h10f == _T_12323 ? mem_271 : _GEN_275;
  assign _GEN_277 = 11'h110 == _T_12323 ? mem_272 : _GEN_276;
  assign _GEN_278 = 11'h111 == _T_12323 ? mem_273 : _GEN_277;
  assign _GEN_279 = 11'h112 == _T_12323 ? mem_274 : _GEN_278;
  assign _GEN_280 = 11'h113 == _T_12323 ? mem_275 : _GEN_279;
  assign _GEN_281 = 11'h114 == _T_12323 ? mem_276 : _GEN_280;
  assign _GEN_282 = 11'h115 == _T_12323 ? mem_277 : _GEN_281;
  assign _GEN_283 = 11'h116 == _T_12323 ? mem_278 : _GEN_282;
  assign _GEN_284 = 11'h117 == _T_12323 ? mem_279 : _GEN_283;
  assign _GEN_285 = 11'h118 == _T_12323 ? mem_280 : _GEN_284;
  assign _GEN_286 = 11'h119 == _T_12323 ? mem_281 : _GEN_285;
  assign _GEN_287 = 11'h11a == _T_12323 ? mem_282 : _GEN_286;
  assign _GEN_288 = 11'h11b == _T_12323 ? mem_283 : _GEN_287;
  assign _GEN_289 = 11'h11c == _T_12323 ? mem_284 : _GEN_288;
  assign _GEN_290 = 11'h11d == _T_12323 ? mem_285 : _GEN_289;
  assign _GEN_291 = 11'h11e == _T_12323 ? mem_286 : _GEN_290;
  assign _GEN_292 = 11'h11f == _T_12323 ? mem_287 : _GEN_291;
  assign _GEN_293 = 11'h120 == _T_12323 ? mem_288 : _GEN_292;
  assign _GEN_294 = 11'h121 == _T_12323 ? mem_289 : _GEN_293;
  assign _GEN_295 = 11'h122 == _T_12323 ? mem_290 : _GEN_294;
  assign _GEN_296 = 11'h123 == _T_12323 ? mem_291 : _GEN_295;
  assign _GEN_297 = 11'h124 == _T_12323 ? mem_292 : _GEN_296;
  assign _GEN_298 = 11'h125 == _T_12323 ? mem_293 : _GEN_297;
  assign _GEN_299 = 11'h126 == _T_12323 ? mem_294 : _GEN_298;
  assign _GEN_300 = 11'h127 == _T_12323 ? mem_295 : _GEN_299;
  assign _GEN_301 = 11'h128 == _T_12323 ? mem_296 : _GEN_300;
  assign _GEN_302 = 11'h129 == _T_12323 ? mem_297 : _GEN_301;
  assign _GEN_303 = 11'h12a == _T_12323 ? mem_298 : _GEN_302;
  assign _GEN_304 = 11'h12b == _T_12323 ? mem_299 : _GEN_303;
  assign _GEN_305 = 11'h12c == _T_12323 ? mem_300 : _GEN_304;
  assign _GEN_306 = 11'h12d == _T_12323 ? mem_301 : _GEN_305;
  assign _GEN_307 = 11'h12e == _T_12323 ? mem_302 : _GEN_306;
  assign _GEN_308 = 11'h12f == _T_12323 ? mem_303 : _GEN_307;
  assign _GEN_309 = 11'h130 == _T_12323 ? mem_304 : _GEN_308;
  assign _GEN_310 = 11'h131 == _T_12323 ? mem_305 : _GEN_309;
  assign _GEN_311 = 11'h132 == _T_12323 ? mem_306 : _GEN_310;
  assign _GEN_312 = 11'h133 == _T_12323 ? mem_307 : _GEN_311;
  assign _GEN_313 = 11'h134 == _T_12323 ? mem_308 : _GEN_312;
  assign _GEN_314 = 11'h135 == _T_12323 ? mem_309 : _GEN_313;
  assign _GEN_315 = 11'h136 == _T_12323 ? mem_310 : _GEN_314;
  assign _GEN_316 = 11'h137 == _T_12323 ? mem_311 : _GEN_315;
  assign _GEN_317 = 11'h138 == _T_12323 ? mem_312 : _GEN_316;
  assign _GEN_318 = 11'h139 == _T_12323 ? mem_313 : _GEN_317;
  assign _GEN_319 = 11'h13a == _T_12323 ? mem_314 : _GEN_318;
  assign _GEN_320 = 11'h13b == _T_12323 ? mem_315 : _GEN_319;
  assign _GEN_321 = 11'h13c == _T_12323 ? mem_316 : _GEN_320;
  assign _GEN_322 = 11'h13d == _T_12323 ? mem_317 : _GEN_321;
  assign _GEN_323 = 11'h13e == _T_12323 ? mem_318 : _GEN_322;
  assign _GEN_324 = 11'h13f == _T_12323 ? mem_319 : _GEN_323;
  assign _GEN_325 = 11'h140 == _T_12323 ? mem_320 : _GEN_324;
  assign _GEN_326 = 11'h141 == _T_12323 ? mem_321 : _GEN_325;
  assign _GEN_327 = 11'h142 == _T_12323 ? mem_322 : _GEN_326;
  assign _GEN_328 = 11'h143 == _T_12323 ? mem_323 : _GEN_327;
  assign _GEN_329 = 11'h144 == _T_12323 ? mem_324 : _GEN_328;
  assign _GEN_330 = 11'h145 == _T_12323 ? mem_325 : _GEN_329;
  assign _GEN_331 = 11'h146 == _T_12323 ? mem_326 : _GEN_330;
  assign _GEN_332 = 11'h147 == _T_12323 ? mem_327 : _GEN_331;
  assign _GEN_333 = 11'h148 == _T_12323 ? mem_328 : _GEN_332;
  assign _GEN_334 = 11'h149 == _T_12323 ? mem_329 : _GEN_333;
  assign _GEN_335 = 11'h14a == _T_12323 ? mem_330 : _GEN_334;
  assign _GEN_336 = 11'h14b == _T_12323 ? mem_331 : _GEN_335;
  assign _GEN_337 = 11'h14c == _T_12323 ? mem_332 : _GEN_336;
  assign _GEN_338 = 11'h14d == _T_12323 ? mem_333 : _GEN_337;
  assign _GEN_339 = 11'h14e == _T_12323 ? mem_334 : _GEN_338;
  assign _GEN_340 = 11'h14f == _T_12323 ? mem_335 : _GEN_339;
  assign _GEN_341 = 11'h150 == _T_12323 ? mem_336 : _GEN_340;
  assign _GEN_342 = 11'h151 == _T_12323 ? mem_337 : _GEN_341;
  assign _GEN_343 = 11'h152 == _T_12323 ? mem_338 : _GEN_342;
  assign _GEN_344 = 11'h153 == _T_12323 ? mem_339 : _GEN_343;
  assign _GEN_345 = 11'h154 == _T_12323 ? mem_340 : _GEN_344;
  assign _GEN_346 = 11'h155 == _T_12323 ? mem_341 : _GEN_345;
  assign _GEN_347 = 11'h156 == _T_12323 ? mem_342 : _GEN_346;
  assign _GEN_348 = 11'h157 == _T_12323 ? mem_343 : _GEN_347;
  assign _GEN_349 = 11'h158 == _T_12323 ? mem_344 : _GEN_348;
  assign _GEN_350 = 11'h159 == _T_12323 ? mem_345 : _GEN_349;
  assign _GEN_351 = 11'h15a == _T_12323 ? mem_346 : _GEN_350;
  assign _GEN_352 = 11'h15b == _T_12323 ? mem_347 : _GEN_351;
  assign _GEN_353 = 11'h15c == _T_12323 ? mem_348 : _GEN_352;
  assign _GEN_354 = 11'h15d == _T_12323 ? mem_349 : _GEN_353;
  assign _GEN_355 = 11'h15e == _T_12323 ? mem_350 : _GEN_354;
  assign _GEN_356 = 11'h15f == _T_12323 ? mem_351 : _GEN_355;
  assign _GEN_357 = 11'h160 == _T_12323 ? mem_352 : _GEN_356;
  assign _GEN_358 = 11'h161 == _T_12323 ? mem_353 : _GEN_357;
  assign _GEN_359 = 11'h162 == _T_12323 ? mem_354 : _GEN_358;
  assign _GEN_360 = 11'h163 == _T_12323 ? mem_355 : _GEN_359;
  assign _GEN_361 = 11'h164 == _T_12323 ? mem_356 : _GEN_360;
  assign _GEN_362 = 11'h165 == _T_12323 ? mem_357 : _GEN_361;
  assign _GEN_363 = 11'h166 == _T_12323 ? mem_358 : _GEN_362;
  assign _GEN_364 = 11'h167 == _T_12323 ? mem_359 : _GEN_363;
  assign _GEN_365 = 11'h168 == _T_12323 ? mem_360 : _GEN_364;
  assign _GEN_366 = 11'h169 == _T_12323 ? mem_361 : _GEN_365;
  assign _GEN_367 = 11'h16a == _T_12323 ? mem_362 : _GEN_366;
  assign _GEN_368 = 11'h16b == _T_12323 ? mem_363 : _GEN_367;
  assign _GEN_369 = 11'h16c == _T_12323 ? mem_364 : _GEN_368;
  assign _GEN_370 = 11'h16d == _T_12323 ? mem_365 : _GEN_369;
  assign _GEN_371 = 11'h16e == _T_12323 ? mem_366 : _GEN_370;
  assign _GEN_372 = 11'h16f == _T_12323 ? mem_367 : _GEN_371;
  assign _GEN_373 = 11'h170 == _T_12323 ? mem_368 : _GEN_372;
  assign _GEN_374 = 11'h171 == _T_12323 ? mem_369 : _GEN_373;
  assign _GEN_375 = 11'h172 == _T_12323 ? mem_370 : _GEN_374;
  assign _GEN_376 = 11'h173 == _T_12323 ? mem_371 : _GEN_375;
  assign _GEN_377 = 11'h174 == _T_12323 ? mem_372 : _GEN_376;
  assign _GEN_378 = 11'h175 == _T_12323 ? mem_373 : _GEN_377;
  assign _GEN_379 = 11'h176 == _T_12323 ? mem_374 : _GEN_378;
  assign _GEN_380 = 11'h177 == _T_12323 ? mem_375 : _GEN_379;
  assign _GEN_381 = 11'h178 == _T_12323 ? mem_376 : _GEN_380;
  assign _GEN_382 = 11'h179 == _T_12323 ? mem_377 : _GEN_381;
  assign _GEN_383 = 11'h17a == _T_12323 ? mem_378 : _GEN_382;
  assign _GEN_384 = 11'h17b == _T_12323 ? mem_379 : _GEN_383;
  assign _GEN_385 = 11'h17c == _T_12323 ? mem_380 : _GEN_384;
  assign _GEN_386 = 11'h17d == _T_12323 ? mem_381 : _GEN_385;
  assign _GEN_387 = 11'h17e == _T_12323 ? mem_382 : _GEN_386;
  assign _GEN_388 = 11'h17f == _T_12323 ? mem_383 : _GEN_387;
  assign _GEN_389 = 11'h180 == _T_12323 ? mem_384 : _GEN_388;
  assign _GEN_390 = 11'h181 == _T_12323 ? mem_385 : _GEN_389;
  assign _GEN_391 = 11'h182 == _T_12323 ? mem_386 : _GEN_390;
  assign _GEN_392 = 11'h183 == _T_12323 ? mem_387 : _GEN_391;
  assign _GEN_393 = 11'h184 == _T_12323 ? mem_388 : _GEN_392;
  assign _GEN_394 = 11'h185 == _T_12323 ? mem_389 : _GEN_393;
  assign _GEN_395 = 11'h186 == _T_12323 ? mem_390 : _GEN_394;
  assign _GEN_396 = 11'h187 == _T_12323 ? mem_391 : _GEN_395;
  assign _GEN_397 = 11'h188 == _T_12323 ? mem_392 : _GEN_396;
  assign _GEN_398 = 11'h189 == _T_12323 ? mem_393 : _GEN_397;
  assign _GEN_399 = 11'h18a == _T_12323 ? mem_394 : _GEN_398;
  assign _GEN_400 = 11'h18b == _T_12323 ? mem_395 : _GEN_399;
  assign _GEN_401 = 11'h18c == _T_12323 ? mem_396 : _GEN_400;
  assign _GEN_402 = 11'h18d == _T_12323 ? mem_397 : _GEN_401;
  assign _GEN_403 = 11'h18e == _T_12323 ? mem_398 : _GEN_402;
  assign _GEN_404 = 11'h18f == _T_12323 ? mem_399 : _GEN_403;
  assign _GEN_405 = 11'h190 == _T_12323 ? mem_400 : _GEN_404;
  assign _GEN_406 = 11'h191 == _T_12323 ? mem_401 : _GEN_405;
  assign _GEN_407 = 11'h192 == _T_12323 ? mem_402 : _GEN_406;
  assign _GEN_408 = 11'h193 == _T_12323 ? mem_403 : _GEN_407;
  assign _GEN_409 = 11'h194 == _T_12323 ? mem_404 : _GEN_408;
  assign _GEN_410 = 11'h195 == _T_12323 ? mem_405 : _GEN_409;
  assign _GEN_411 = 11'h196 == _T_12323 ? mem_406 : _GEN_410;
  assign _GEN_412 = 11'h197 == _T_12323 ? mem_407 : _GEN_411;
  assign _GEN_413 = 11'h198 == _T_12323 ? mem_408 : _GEN_412;
  assign _GEN_414 = 11'h199 == _T_12323 ? mem_409 : _GEN_413;
  assign _GEN_415 = 11'h19a == _T_12323 ? mem_410 : _GEN_414;
  assign _GEN_416 = 11'h19b == _T_12323 ? mem_411 : _GEN_415;
  assign _GEN_417 = 11'h19c == _T_12323 ? mem_412 : _GEN_416;
  assign _GEN_418 = 11'h19d == _T_12323 ? mem_413 : _GEN_417;
  assign _GEN_419 = 11'h19e == _T_12323 ? mem_414 : _GEN_418;
  assign _GEN_420 = 11'h19f == _T_12323 ? mem_415 : _GEN_419;
  assign _GEN_421 = 11'h1a0 == _T_12323 ? mem_416 : _GEN_420;
  assign _GEN_422 = 11'h1a1 == _T_12323 ? mem_417 : _GEN_421;
  assign _GEN_423 = 11'h1a2 == _T_12323 ? mem_418 : _GEN_422;
  assign _GEN_424 = 11'h1a3 == _T_12323 ? mem_419 : _GEN_423;
  assign _GEN_425 = 11'h1a4 == _T_12323 ? mem_420 : _GEN_424;
  assign _GEN_426 = 11'h1a5 == _T_12323 ? mem_421 : _GEN_425;
  assign _GEN_427 = 11'h1a6 == _T_12323 ? mem_422 : _GEN_426;
  assign _GEN_428 = 11'h1a7 == _T_12323 ? mem_423 : _GEN_427;
  assign _GEN_429 = 11'h1a8 == _T_12323 ? mem_424 : _GEN_428;
  assign _GEN_430 = 11'h1a9 == _T_12323 ? mem_425 : _GEN_429;
  assign _GEN_431 = 11'h1aa == _T_12323 ? mem_426 : _GEN_430;
  assign _GEN_432 = 11'h1ab == _T_12323 ? mem_427 : _GEN_431;
  assign _GEN_433 = 11'h1ac == _T_12323 ? mem_428 : _GEN_432;
  assign _GEN_434 = 11'h1ad == _T_12323 ? mem_429 : _GEN_433;
  assign _GEN_435 = 11'h1ae == _T_12323 ? mem_430 : _GEN_434;
  assign _GEN_436 = 11'h1af == _T_12323 ? mem_431 : _GEN_435;
  assign _GEN_437 = 11'h1b0 == _T_12323 ? mem_432 : _GEN_436;
  assign _GEN_438 = 11'h1b1 == _T_12323 ? mem_433 : _GEN_437;
  assign _GEN_439 = 11'h1b2 == _T_12323 ? mem_434 : _GEN_438;
  assign _GEN_440 = 11'h1b3 == _T_12323 ? mem_435 : _GEN_439;
  assign _GEN_441 = 11'h1b4 == _T_12323 ? mem_436 : _GEN_440;
  assign _GEN_442 = 11'h1b5 == _T_12323 ? mem_437 : _GEN_441;
  assign _GEN_443 = 11'h1b6 == _T_12323 ? mem_438 : _GEN_442;
  assign _GEN_444 = 11'h1b7 == _T_12323 ? mem_439 : _GEN_443;
  assign _GEN_445 = 11'h1b8 == _T_12323 ? mem_440 : _GEN_444;
  assign _GEN_446 = 11'h1b9 == _T_12323 ? mem_441 : _GEN_445;
  assign _GEN_447 = 11'h1ba == _T_12323 ? mem_442 : _GEN_446;
  assign _GEN_448 = 11'h1bb == _T_12323 ? mem_443 : _GEN_447;
  assign _GEN_449 = 11'h1bc == _T_12323 ? mem_444 : _GEN_448;
  assign _GEN_450 = 11'h1bd == _T_12323 ? mem_445 : _GEN_449;
  assign _GEN_451 = 11'h1be == _T_12323 ? mem_446 : _GEN_450;
  assign _GEN_452 = 11'h1bf == _T_12323 ? mem_447 : _GEN_451;
  assign _GEN_453 = 11'h1c0 == _T_12323 ? mem_448 : _GEN_452;
  assign _GEN_454 = 11'h1c1 == _T_12323 ? mem_449 : _GEN_453;
  assign _GEN_455 = 11'h1c2 == _T_12323 ? mem_450 : _GEN_454;
  assign _GEN_456 = 11'h1c3 == _T_12323 ? mem_451 : _GEN_455;
  assign _GEN_457 = 11'h1c4 == _T_12323 ? mem_452 : _GEN_456;
  assign _GEN_458 = 11'h1c5 == _T_12323 ? mem_453 : _GEN_457;
  assign _GEN_459 = 11'h1c6 == _T_12323 ? mem_454 : _GEN_458;
  assign _GEN_460 = 11'h1c7 == _T_12323 ? mem_455 : _GEN_459;
  assign _GEN_461 = 11'h1c8 == _T_12323 ? mem_456 : _GEN_460;
  assign _GEN_462 = 11'h1c9 == _T_12323 ? mem_457 : _GEN_461;
  assign _GEN_463 = 11'h1ca == _T_12323 ? mem_458 : _GEN_462;
  assign _GEN_464 = 11'h1cb == _T_12323 ? mem_459 : _GEN_463;
  assign _GEN_465 = 11'h1cc == _T_12323 ? mem_460 : _GEN_464;
  assign _GEN_466 = 11'h1cd == _T_12323 ? mem_461 : _GEN_465;
  assign _GEN_467 = 11'h1ce == _T_12323 ? mem_462 : _GEN_466;
  assign _GEN_468 = 11'h1cf == _T_12323 ? mem_463 : _GEN_467;
  assign _GEN_469 = 11'h1d0 == _T_12323 ? mem_464 : _GEN_468;
  assign _GEN_470 = 11'h1d1 == _T_12323 ? mem_465 : _GEN_469;
  assign _GEN_471 = 11'h1d2 == _T_12323 ? mem_466 : _GEN_470;
  assign _GEN_472 = 11'h1d3 == _T_12323 ? mem_467 : _GEN_471;
  assign _GEN_473 = 11'h1d4 == _T_12323 ? mem_468 : _GEN_472;
  assign _GEN_474 = 11'h1d5 == _T_12323 ? mem_469 : _GEN_473;
  assign _GEN_475 = 11'h1d6 == _T_12323 ? mem_470 : _GEN_474;
  assign _GEN_476 = 11'h1d7 == _T_12323 ? mem_471 : _GEN_475;
  assign _GEN_477 = 11'h1d8 == _T_12323 ? mem_472 : _GEN_476;
  assign _GEN_478 = 11'h1d9 == _T_12323 ? mem_473 : _GEN_477;
  assign _GEN_479 = 11'h1da == _T_12323 ? mem_474 : _GEN_478;
  assign _GEN_480 = 11'h1db == _T_12323 ? mem_475 : _GEN_479;
  assign _GEN_481 = 11'h1dc == _T_12323 ? mem_476 : _GEN_480;
  assign _GEN_482 = 11'h1dd == _T_12323 ? mem_477 : _GEN_481;
  assign _GEN_483 = 11'h1de == _T_12323 ? mem_478 : _GEN_482;
  assign _GEN_484 = 11'h1df == _T_12323 ? mem_479 : _GEN_483;
  assign _GEN_485 = 11'h1e0 == _T_12323 ? mem_480 : _GEN_484;
  assign _GEN_486 = 11'h1e1 == _T_12323 ? mem_481 : _GEN_485;
  assign _GEN_487 = 11'h1e2 == _T_12323 ? mem_482 : _GEN_486;
  assign _GEN_488 = 11'h1e3 == _T_12323 ? mem_483 : _GEN_487;
  assign _GEN_489 = 11'h1e4 == _T_12323 ? mem_484 : _GEN_488;
  assign _GEN_490 = 11'h1e5 == _T_12323 ? mem_485 : _GEN_489;
  assign _GEN_491 = 11'h1e6 == _T_12323 ? mem_486 : _GEN_490;
  assign _GEN_492 = 11'h1e7 == _T_12323 ? mem_487 : _GEN_491;
  assign _GEN_493 = 11'h1e8 == _T_12323 ? mem_488 : _GEN_492;
  assign _GEN_494 = 11'h1e9 == _T_12323 ? mem_489 : _GEN_493;
  assign _GEN_495 = 11'h1ea == _T_12323 ? mem_490 : _GEN_494;
  assign _GEN_496 = 11'h1eb == _T_12323 ? mem_491 : _GEN_495;
  assign _GEN_497 = 11'h1ec == _T_12323 ? mem_492 : _GEN_496;
  assign _GEN_498 = 11'h1ed == _T_12323 ? mem_493 : _GEN_497;
  assign _GEN_499 = 11'h1ee == _T_12323 ? mem_494 : _GEN_498;
  assign _GEN_500 = 11'h1ef == _T_12323 ? mem_495 : _GEN_499;
  assign _GEN_501 = 11'h1f0 == _T_12323 ? mem_496 : _GEN_500;
  assign _GEN_502 = 11'h1f1 == _T_12323 ? mem_497 : _GEN_501;
  assign _GEN_503 = 11'h1f2 == _T_12323 ? mem_498 : _GEN_502;
  assign _GEN_504 = 11'h1f3 == _T_12323 ? mem_499 : _GEN_503;
  assign _GEN_505 = 11'h1f4 == _T_12323 ? mem_500 : _GEN_504;
  assign _GEN_506 = 11'h1f5 == _T_12323 ? mem_501 : _GEN_505;
  assign _GEN_507 = 11'h1f6 == _T_12323 ? mem_502 : _GEN_506;
  assign _GEN_508 = 11'h1f7 == _T_12323 ? mem_503 : _GEN_507;
  assign _GEN_509 = 11'h1f8 == _T_12323 ? mem_504 : _GEN_508;
  assign _GEN_510 = 11'h1f9 == _T_12323 ? mem_505 : _GEN_509;
  assign _GEN_511 = 11'h1fa == _T_12323 ? mem_506 : _GEN_510;
  assign _GEN_512 = 11'h1fb == _T_12323 ? mem_507 : _GEN_511;
  assign _GEN_513 = 11'h1fc == _T_12323 ? mem_508 : _GEN_512;
  assign _GEN_514 = 11'h1fd == _T_12323 ? mem_509 : _GEN_513;
  assign _GEN_515 = 11'h1fe == _T_12323 ? mem_510 : _GEN_514;
  assign _GEN_516 = 11'h1ff == _T_12323 ? mem_511 : _GEN_515;
  assign _GEN_517 = 11'h200 == _T_12323 ? mem_512 : _GEN_516;
  assign _GEN_518 = 11'h201 == _T_12323 ? mem_513 : _GEN_517;
  assign _GEN_519 = 11'h202 == _T_12323 ? mem_514 : _GEN_518;
  assign _GEN_520 = 11'h203 == _T_12323 ? mem_515 : _GEN_519;
  assign _GEN_521 = 11'h204 == _T_12323 ? mem_516 : _GEN_520;
  assign _GEN_522 = 11'h205 == _T_12323 ? mem_517 : _GEN_521;
  assign _GEN_523 = 11'h206 == _T_12323 ? mem_518 : _GEN_522;
  assign _GEN_524 = 11'h207 == _T_12323 ? mem_519 : _GEN_523;
  assign _GEN_525 = 11'h208 == _T_12323 ? mem_520 : _GEN_524;
  assign _GEN_526 = 11'h209 == _T_12323 ? mem_521 : _GEN_525;
  assign _GEN_527 = 11'h20a == _T_12323 ? mem_522 : _GEN_526;
  assign _GEN_528 = 11'h20b == _T_12323 ? mem_523 : _GEN_527;
  assign _GEN_529 = 11'h20c == _T_12323 ? mem_524 : _GEN_528;
  assign _GEN_530 = 11'h20d == _T_12323 ? mem_525 : _GEN_529;
  assign _GEN_531 = 11'h20e == _T_12323 ? mem_526 : _GEN_530;
  assign _GEN_532 = 11'h20f == _T_12323 ? mem_527 : _GEN_531;
  assign _GEN_533 = 11'h210 == _T_12323 ? mem_528 : _GEN_532;
  assign _GEN_534 = 11'h211 == _T_12323 ? mem_529 : _GEN_533;
  assign _GEN_535 = 11'h212 == _T_12323 ? mem_530 : _GEN_534;
  assign _GEN_536 = 11'h213 == _T_12323 ? mem_531 : _GEN_535;
  assign _GEN_537 = 11'h214 == _T_12323 ? mem_532 : _GEN_536;
  assign _GEN_538 = 11'h215 == _T_12323 ? mem_533 : _GEN_537;
  assign _GEN_539 = 11'h216 == _T_12323 ? mem_534 : _GEN_538;
  assign _GEN_540 = 11'h217 == _T_12323 ? mem_535 : _GEN_539;
  assign _GEN_541 = 11'h218 == _T_12323 ? mem_536 : _GEN_540;
  assign _GEN_542 = 11'h219 == _T_12323 ? mem_537 : _GEN_541;
  assign _GEN_543 = 11'h21a == _T_12323 ? mem_538 : _GEN_542;
  assign _GEN_544 = 11'h21b == _T_12323 ? mem_539 : _GEN_543;
  assign _GEN_545 = 11'h21c == _T_12323 ? mem_540 : _GEN_544;
  assign _GEN_546 = 11'h21d == _T_12323 ? mem_541 : _GEN_545;
  assign _GEN_547 = 11'h21e == _T_12323 ? mem_542 : _GEN_546;
  assign _GEN_548 = 11'h21f == _T_12323 ? mem_543 : _GEN_547;
  assign _GEN_549 = 11'h220 == _T_12323 ? mem_544 : _GEN_548;
  assign _GEN_550 = 11'h221 == _T_12323 ? mem_545 : _GEN_549;
  assign _GEN_551 = 11'h222 == _T_12323 ? mem_546 : _GEN_550;
  assign _GEN_552 = 11'h223 == _T_12323 ? mem_547 : _GEN_551;
  assign _GEN_553 = 11'h224 == _T_12323 ? mem_548 : _GEN_552;
  assign _GEN_554 = 11'h225 == _T_12323 ? mem_549 : _GEN_553;
  assign _GEN_555 = 11'h226 == _T_12323 ? mem_550 : _GEN_554;
  assign _GEN_556 = 11'h227 == _T_12323 ? mem_551 : _GEN_555;
  assign _GEN_557 = 11'h228 == _T_12323 ? mem_552 : _GEN_556;
  assign _GEN_558 = 11'h229 == _T_12323 ? mem_553 : _GEN_557;
  assign _GEN_559 = 11'h22a == _T_12323 ? mem_554 : _GEN_558;
  assign _GEN_560 = 11'h22b == _T_12323 ? mem_555 : _GEN_559;
  assign _GEN_561 = 11'h22c == _T_12323 ? mem_556 : _GEN_560;
  assign _GEN_562 = 11'h22d == _T_12323 ? mem_557 : _GEN_561;
  assign _GEN_563 = 11'h22e == _T_12323 ? mem_558 : _GEN_562;
  assign _GEN_564 = 11'h22f == _T_12323 ? mem_559 : _GEN_563;
  assign _GEN_565 = 11'h230 == _T_12323 ? mem_560 : _GEN_564;
  assign _GEN_566 = 11'h231 == _T_12323 ? mem_561 : _GEN_565;
  assign _GEN_567 = 11'h232 == _T_12323 ? mem_562 : _GEN_566;
  assign _GEN_568 = 11'h233 == _T_12323 ? mem_563 : _GEN_567;
  assign _GEN_569 = 11'h234 == _T_12323 ? mem_564 : _GEN_568;
  assign _GEN_570 = 11'h235 == _T_12323 ? mem_565 : _GEN_569;
  assign _GEN_571 = 11'h236 == _T_12323 ? mem_566 : _GEN_570;
  assign _GEN_572 = 11'h237 == _T_12323 ? mem_567 : _GEN_571;
  assign _GEN_573 = 11'h238 == _T_12323 ? mem_568 : _GEN_572;
  assign _GEN_574 = 11'h239 == _T_12323 ? mem_569 : _GEN_573;
  assign _GEN_575 = 11'h23a == _T_12323 ? mem_570 : _GEN_574;
  assign _GEN_576 = 11'h23b == _T_12323 ? mem_571 : _GEN_575;
  assign _GEN_577 = 11'h23c == _T_12323 ? mem_572 : _GEN_576;
  assign _GEN_578 = 11'h23d == _T_12323 ? mem_573 : _GEN_577;
  assign _GEN_579 = 11'h23e == _T_12323 ? mem_574 : _GEN_578;
  assign _GEN_580 = 11'h23f == _T_12323 ? mem_575 : _GEN_579;
  assign _GEN_581 = 11'h240 == _T_12323 ? mem_576 : _GEN_580;
  assign _GEN_582 = 11'h241 == _T_12323 ? mem_577 : _GEN_581;
  assign _GEN_583 = 11'h242 == _T_12323 ? mem_578 : _GEN_582;
  assign _GEN_584 = 11'h243 == _T_12323 ? mem_579 : _GEN_583;
  assign _GEN_585 = 11'h244 == _T_12323 ? mem_580 : _GEN_584;
  assign _GEN_586 = 11'h245 == _T_12323 ? mem_581 : _GEN_585;
  assign _GEN_587 = 11'h246 == _T_12323 ? mem_582 : _GEN_586;
  assign _GEN_588 = 11'h247 == _T_12323 ? mem_583 : _GEN_587;
  assign _GEN_589 = 11'h248 == _T_12323 ? mem_584 : _GEN_588;
  assign _GEN_590 = 11'h249 == _T_12323 ? mem_585 : _GEN_589;
  assign _GEN_591 = 11'h24a == _T_12323 ? mem_586 : _GEN_590;
  assign _GEN_592 = 11'h24b == _T_12323 ? mem_587 : _GEN_591;
  assign _GEN_593 = 11'h24c == _T_12323 ? mem_588 : _GEN_592;
  assign _GEN_594 = 11'h24d == _T_12323 ? mem_589 : _GEN_593;
  assign _GEN_595 = 11'h24e == _T_12323 ? mem_590 : _GEN_594;
  assign _GEN_596 = 11'h24f == _T_12323 ? mem_591 : _GEN_595;
  assign _GEN_597 = 11'h250 == _T_12323 ? mem_592 : _GEN_596;
  assign _GEN_598 = 11'h251 == _T_12323 ? mem_593 : _GEN_597;
  assign _GEN_599 = 11'h252 == _T_12323 ? mem_594 : _GEN_598;
  assign _GEN_600 = 11'h253 == _T_12323 ? mem_595 : _GEN_599;
  assign _GEN_601 = 11'h254 == _T_12323 ? mem_596 : _GEN_600;
  assign _GEN_602 = 11'h255 == _T_12323 ? mem_597 : _GEN_601;
  assign _GEN_603 = 11'h256 == _T_12323 ? mem_598 : _GEN_602;
  assign _GEN_604 = 11'h257 == _T_12323 ? mem_599 : _GEN_603;
  assign _GEN_605 = 11'h258 == _T_12323 ? mem_600 : _GEN_604;
  assign _GEN_606 = 11'h259 == _T_12323 ? mem_601 : _GEN_605;
  assign _GEN_607 = 11'h25a == _T_12323 ? mem_602 : _GEN_606;
  assign _GEN_608 = 11'h25b == _T_12323 ? mem_603 : _GEN_607;
  assign _GEN_609 = 11'h25c == _T_12323 ? mem_604 : _GEN_608;
  assign _GEN_610 = 11'h25d == _T_12323 ? mem_605 : _GEN_609;
  assign _GEN_611 = 11'h25e == _T_12323 ? mem_606 : _GEN_610;
  assign _GEN_612 = 11'h25f == _T_12323 ? mem_607 : _GEN_611;
  assign _GEN_613 = 11'h260 == _T_12323 ? mem_608 : _GEN_612;
  assign _GEN_614 = 11'h261 == _T_12323 ? mem_609 : _GEN_613;
  assign _GEN_615 = 11'h262 == _T_12323 ? mem_610 : _GEN_614;
  assign _GEN_616 = 11'h263 == _T_12323 ? mem_611 : _GEN_615;
  assign _GEN_617 = 11'h264 == _T_12323 ? mem_612 : _GEN_616;
  assign _GEN_618 = 11'h265 == _T_12323 ? mem_613 : _GEN_617;
  assign _GEN_619 = 11'h266 == _T_12323 ? mem_614 : _GEN_618;
  assign _GEN_620 = 11'h267 == _T_12323 ? mem_615 : _GEN_619;
  assign _GEN_621 = 11'h268 == _T_12323 ? mem_616 : _GEN_620;
  assign _GEN_622 = 11'h269 == _T_12323 ? mem_617 : _GEN_621;
  assign _GEN_623 = 11'h26a == _T_12323 ? mem_618 : _GEN_622;
  assign _GEN_624 = 11'h26b == _T_12323 ? mem_619 : _GEN_623;
  assign _GEN_625 = 11'h26c == _T_12323 ? mem_620 : _GEN_624;
  assign _GEN_626 = 11'h26d == _T_12323 ? mem_621 : _GEN_625;
  assign _GEN_627 = 11'h26e == _T_12323 ? mem_622 : _GEN_626;
  assign _GEN_628 = 11'h26f == _T_12323 ? mem_623 : _GEN_627;
  assign _GEN_629 = 11'h270 == _T_12323 ? mem_624 : _GEN_628;
  assign _GEN_630 = 11'h271 == _T_12323 ? mem_625 : _GEN_629;
  assign _GEN_631 = 11'h272 == _T_12323 ? mem_626 : _GEN_630;
  assign _GEN_632 = 11'h273 == _T_12323 ? mem_627 : _GEN_631;
  assign _GEN_633 = 11'h274 == _T_12323 ? mem_628 : _GEN_632;
  assign _GEN_634 = 11'h275 == _T_12323 ? mem_629 : _GEN_633;
  assign _GEN_635 = 11'h276 == _T_12323 ? mem_630 : _GEN_634;
  assign _GEN_636 = 11'h277 == _T_12323 ? mem_631 : _GEN_635;
  assign _GEN_637 = 11'h278 == _T_12323 ? mem_632 : _GEN_636;
  assign _GEN_638 = 11'h279 == _T_12323 ? mem_633 : _GEN_637;
  assign _GEN_639 = 11'h27a == _T_12323 ? mem_634 : _GEN_638;
  assign _GEN_640 = 11'h27b == _T_12323 ? mem_635 : _GEN_639;
  assign _GEN_641 = 11'h27c == _T_12323 ? mem_636 : _GEN_640;
  assign _GEN_642 = 11'h27d == _T_12323 ? mem_637 : _GEN_641;
  assign _GEN_643 = 11'h27e == _T_12323 ? mem_638 : _GEN_642;
  assign _GEN_644 = 11'h27f == _T_12323 ? mem_639 : _GEN_643;
  assign _GEN_645 = 11'h280 == _T_12323 ? mem_640 : _GEN_644;
  assign _GEN_646 = 11'h281 == _T_12323 ? mem_641 : _GEN_645;
  assign _GEN_647 = 11'h282 == _T_12323 ? mem_642 : _GEN_646;
  assign _GEN_648 = 11'h283 == _T_12323 ? mem_643 : _GEN_647;
  assign _GEN_649 = 11'h284 == _T_12323 ? mem_644 : _GEN_648;
  assign _GEN_650 = 11'h285 == _T_12323 ? mem_645 : _GEN_649;
  assign _GEN_651 = 11'h286 == _T_12323 ? mem_646 : _GEN_650;
  assign _GEN_652 = 11'h287 == _T_12323 ? mem_647 : _GEN_651;
  assign _GEN_653 = 11'h288 == _T_12323 ? mem_648 : _GEN_652;
  assign _GEN_654 = 11'h289 == _T_12323 ? mem_649 : _GEN_653;
  assign _GEN_655 = 11'h28a == _T_12323 ? mem_650 : _GEN_654;
  assign _GEN_656 = 11'h28b == _T_12323 ? mem_651 : _GEN_655;
  assign _GEN_657 = 11'h28c == _T_12323 ? mem_652 : _GEN_656;
  assign _GEN_658 = 11'h28d == _T_12323 ? mem_653 : _GEN_657;
  assign _GEN_659 = 11'h28e == _T_12323 ? mem_654 : _GEN_658;
  assign _GEN_660 = 11'h28f == _T_12323 ? mem_655 : _GEN_659;
  assign _GEN_661 = 11'h290 == _T_12323 ? mem_656 : _GEN_660;
  assign _GEN_662 = 11'h291 == _T_12323 ? mem_657 : _GEN_661;
  assign _GEN_663 = 11'h292 == _T_12323 ? mem_658 : _GEN_662;
  assign _GEN_664 = 11'h293 == _T_12323 ? mem_659 : _GEN_663;
  assign _GEN_665 = 11'h294 == _T_12323 ? mem_660 : _GEN_664;
  assign _GEN_666 = 11'h295 == _T_12323 ? mem_661 : _GEN_665;
  assign _GEN_667 = 11'h296 == _T_12323 ? mem_662 : _GEN_666;
  assign _GEN_668 = 11'h297 == _T_12323 ? mem_663 : _GEN_667;
  assign _GEN_669 = 11'h298 == _T_12323 ? mem_664 : _GEN_668;
  assign _GEN_670 = 11'h299 == _T_12323 ? mem_665 : _GEN_669;
  assign _GEN_671 = 11'h29a == _T_12323 ? mem_666 : _GEN_670;
  assign _GEN_672 = 11'h29b == _T_12323 ? mem_667 : _GEN_671;
  assign _GEN_673 = 11'h29c == _T_12323 ? mem_668 : _GEN_672;
  assign _GEN_674 = 11'h29d == _T_12323 ? mem_669 : _GEN_673;
  assign _GEN_675 = 11'h29e == _T_12323 ? mem_670 : _GEN_674;
  assign _GEN_676 = 11'h29f == _T_12323 ? mem_671 : _GEN_675;
  assign _GEN_677 = 11'h2a0 == _T_12323 ? mem_672 : _GEN_676;
  assign _GEN_678 = 11'h2a1 == _T_12323 ? mem_673 : _GEN_677;
  assign _GEN_679 = 11'h2a2 == _T_12323 ? mem_674 : _GEN_678;
  assign _GEN_680 = 11'h2a3 == _T_12323 ? mem_675 : _GEN_679;
  assign _GEN_681 = 11'h2a4 == _T_12323 ? mem_676 : _GEN_680;
  assign _GEN_682 = 11'h2a5 == _T_12323 ? mem_677 : _GEN_681;
  assign _GEN_683 = 11'h2a6 == _T_12323 ? mem_678 : _GEN_682;
  assign _GEN_684 = 11'h2a7 == _T_12323 ? mem_679 : _GEN_683;
  assign _GEN_685 = 11'h2a8 == _T_12323 ? mem_680 : _GEN_684;
  assign _GEN_686 = 11'h2a9 == _T_12323 ? mem_681 : _GEN_685;
  assign _GEN_687 = 11'h2aa == _T_12323 ? mem_682 : _GEN_686;
  assign _GEN_688 = 11'h2ab == _T_12323 ? mem_683 : _GEN_687;
  assign _GEN_689 = 11'h2ac == _T_12323 ? mem_684 : _GEN_688;
  assign _GEN_690 = 11'h2ad == _T_12323 ? mem_685 : _GEN_689;
  assign _GEN_691 = 11'h2ae == _T_12323 ? mem_686 : _GEN_690;
  assign _GEN_692 = 11'h2af == _T_12323 ? mem_687 : _GEN_691;
  assign _GEN_693 = 11'h2b0 == _T_12323 ? mem_688 : _GEN_692;
  assign _GEN_694 = 11'h2b1 == _T_12323 ? mem_689 : _GEN_693;
  assign _GEN_695 = 11'h2b2 == _T_12323 ? mem_690 : _GEN_694;
  assign _GEN_696 = 11'h2b3 == _T_12323 ? mem_691 : _GEN_695;
  assign _GEN_697 = 11'h2b4 == _T_12323 ? mem_692 : _GEN_696;
  assign _GEN_698 = 11'h2b5 == _T_12323 ? mem_693 : _GEN_697;
  assign _GEN_699 = 11'h2b6 == _T_12323 ? mem_694 : _GEN_698;
  assign _GEN_700 = 11'h2b7 == _T_12323 ? mem_695 : _GEN_699;
  assign _GEN_701 = 11'h2b8 == _T_12323 ? mem_696 : _GEN_700;
  assign _GEN_702 = 11'h2b9 == _T_12323 ? mem_697 : _GEN_701;
  assign _GEN_703 = 11'h2ba == _T_12323 ? mem_698 : _GEN_702;
  assign _GEN_704 = 11'h2bb == _T_12323 ? mem_699 : _GEN_703;
  assign _GEN_705 = 11'h2bc == _T_12323 ? mem_700 : _GEN_704;
  assign _GEN_706 = 11'h2bd == _T_12323 ? mem_701 : _GEN_705;
  assign _GEN_707 = 11'h2be == _T_12323 ? mem_702 : _GEN_706;
  assign _GEN_708 = 11'h2bf == _T_12323 ? mem_703 : _GEN_707;
  assign _GEN_709 = 11'h2c0 == _T_12323 ? mem_704 : _GEN_708;
  assign _GEN_710 = 11'h2c1 == _T_12323 ? mem_705 : _GEN_709;
  assign _GEN_711 = 11'h2c2 == _T_12323 ? mem_706 : _GEN_710;
  assign _GEN_712 = 11'h2c3 == _T_12323 ? mem_707 : _GEN_711;
  assign _GEN_713 = 11'h2c4 == _T_12323 ? mem_708 : _GEN_712;
  assign _GEN_714 = 11'h2c5 == _T_12323 ? mem_709 : _GEN_713;
  assign _GEN_715 = 11'h2c6 == _T_12323 ? mem_710 : _GEN_714;
  assign _GEN_716 = 11'h2c7 == _T_12323 ? mem_711 : _GEN_715;
  assign _GEN_717 = 11'h2c8 == _T_12323 ? mem_712 : _GEN_716;
  assign _GEN_718 = 11'h2c9 == _T_12323 ? mem_713 : _GEN_717;
  assign _GEN_719 = 11'h2ca == _T_12323 ? mem_714 : _GEN_718;
  assign _GEN_720 = 11'h2cb == _T_12323 ? mem_715 : _GEN_719;
  assign _GEN_721 = 11'h2cc == _T_12323 ? mem_716 : _GEN_720;
  assign _GEN_722 = 11'h2cd == _T_12323 ? mem_717 : _GEN_721;
  assign _GEN_723 = 11'h2ce == _T_12323 ? mem_718 : _GEN_722;
  assign _GEN_724 = 11'h2cf == _T_12323 ? mem_719 : _GEN_723;
  assign _GEN_725 = 11'h2d0 == _T_12323 ? mem_720 : _GEN_724;
  assign _GEN_726 = 11'h2d1 == _T_12323 ? mem_721 : _GEN_725;
  assign _GEN_727 = 11'h2d2 == _T_12323 ? mem_722 : _GEN_726;
  assign _GEN_728 = 11'h2d3 == _T_12323 ? mem_723 : _GEN_727;
  assign _GEN_729 = 11'h2d4 == _T_12323 ? mem_724 : _GEN_728;
  assign _GEN_730 = 11'h2d5 == _T_12323 ? mem_725 : _GEN_729;
  assign _GEN_731 = 11'h2d6 == _T_12323 ? mem_726 : _GEN_730;
  assign _GEN_732 = 11'h2d7 == _T_12323 ? mem_727 : _GEN_731;
  assign _GEN_733 = 11'h2d8 == _T_12323 ? mem_728 : _GEN_732;
  assign _GEN_734 = 11'h2d9 == _T_12323 ? mem_729 : _GEN_733;
  assign _GEN_735 = 11'h2da == _T_12323 ? mem_730 : _GEN_734;
  assign _GEN_736 = 11'h2db == _T_12323 ? mem_731 : _GEN_735;
  assign _GEN_737 = 11'h2dc == _T_12323 ? mem_732 : _GEN_736;
  assign _GEN_738 = 11'h2dd == _T_12323 ? mem_733 : _GEN_737;
  assign _GEN_739 = 11'h2de == _T_12323 ? mem_734 : _GEN_738;
  assign _GEN_740 = 11'h2df == _T_12323 ? mem_735 : _GEN_739;
  assign _GEN_741 = 11'h2e0 == _T_12323 ? mem_736 : _GEN_740;
  assign _GEN_742 = 11'h2e1 == _T_12323 ? mem_737 : _GEN_741;
  assign _GEN_743 = 11'h2e2 == _T_12323 ? mem_738 : _GEN_742;
  assign _GEN_744 = 11'h2e3 == _T_12323 ? mem_739 : _GEN_743;
  assign _GEN_745 = 11'h2e4 == _T_12323 ? mem_740 : _GEN_744;
  assign _GEN_746 = 11'h2e5 == _T_12323 ? mem_741 : _GEN_745;
  assign _GEN_747 = 11'h2e6 == _T_12323 ? mem_742 : _GEN_746;
  assign _GEN_748 = 11'h2e7 == _T_12323 ? mem_743 : _GEN_747;
  assign _GEN_749 = 11'h2e8 == _T_12323 ? mem_744 : _GEN_748;
  assign _GEN_750 = 11'h2e9 == _T_12323 ? mem_745 : _GEN_749;
  assign _GEN_751 = 11'h2ea == _T_12323 ? mem_746 : _GEN_750;
  assign _GEN_752 = 11'h2eb == _T_12323 ? mem_747 : _GEN_751;
  assign _GEN_753 = 11'h2ec == _T_12323 ? mem_748 : _GEN_752;
  assign _GEN_754 = 11'h2ed == _T_12323 ? mem_749 : _GEN_753;
  assign _GEN_755 = 11'h2ee == _T_12323 ? mem_750 : _GEN_754;
  assign _GEN_756 = 11'h2ef == _T_12323 ? mem_751 : _GEN_755;
  assign _GEN_757 = 11'h2f0 == _T_12323 ? mem_752 : _GEN_756;
  assign _GEN_758 = 11'h2f1 == _T_12323 ? mem_753 : _GEN_757;
  assign _GEN_759 = 11'h2f2 == _T_12323 ? mem_754 : _GEN_758;
  assign _GEN_760 = 11'h2f3 == _T_12323 ? mem_755 : _GEN_759;
  assign _GEN_761 = 11'h2f4 == _T_12323 ? mem_756 : _GEN_760;
  assign _GEN_762 = 11'h2f5 == _T_12323 ? mem_757 : _GEN_761;
  assign _GEN_763 = 11'h2f6 == _T_12323 ? mem_758 : _GEN_762;
  assign _GEN_764 = 11'h2f7 == _T_12323 ? mem_759 : _GEN_763;
  assign _GEN_765 = 11'h2f8 == _T_12323 ? mem_760 : _GEN_764;
  assign _GEN_766 = 11'h2f9 == _T_12323 ? mem_761 : _GEN_765;
  assign _GEN_767 = 11'h2fa == _T_12323 ? mem_762 : _GEN_766;
  assign _GEN_768 = 11'h2fb == _T_12323 ? mem_763 : _GEN_767;
  assign _GEN_769 = 11'h2fc == _T_12323 ? mem_764 : _GEN_768;
  assign _GEN_770 = 11'h2fd == _T_12323 ? mem_765 : _GEN_769;
  assign _GEN_771 = 11'h2fe == _T_12323 ? mem_766 : _GEN_770;
  assign _GEN_772 = 11'h2ff == _T_12323 ? mem_767 : _GEN_771;
  assign _GEN_773 = 11'h300 == _T_12323 ? mem_768 : _GEN_772;
  assign _GEN_774 = 11'h301 == _T_12323 ? mem_769 : _GEN_773;
  assign _GEN_775 = 11'h302 == _T_12323 ? mem_770 : _GEN_774;
  assign _GEN_776 = 11'h303 == _T_12323 ? mem_771 : _GEN_775;
  assign _GEN_777 = 11'h304 == _T_12323 ? mem_772 : _GEN_776;
  assign _GEN_778 = 11'h305 == _T_12323 ? mem_773 : _GEN_777;
  assign _GEN_779 = 11'h306 == _T_12323 ? mem_774 : _GEN_778;
  assign _GEN_780 = 11'h307 == _T_12323 ? mem_775 : _GEN_779;
  assign _GEN_781 = 11'h308 == _T_12323 ? mem_776 : _GEN_780;
  assign _GEN_782 = 11'h309 == _T_12323 ? mem_777 : _GEN_781;
  assign _GEN_783 = 11'h30a == _T_12323 ? mem_778 : _GEN_782;
  assign _GEN_784 = 11'h30b == _T_12323 ? mem_779 : _GEN_783;
  assign _GEN_785 = 11'h30c == _T_12323 ? mem_780 : _GEN_784;
  assign _GEN_786 = 11'h30d == _T_12323 ? mem_781 : _GEN_785;
  assign _GEN_787 = 11'h30e == _T_12323 ? mem_782 : _GEN_786;
  assign _GEN_788 = 11'h30f == _T_12323 ? mem_783 : _GEN_787;
  assign _GEN_789 = 11'h310 == _T_12323 ? mem_784 : _GEN_788;
  assign _GEN_790 = 11'h311 == _T_12323 ? mem_785 : _GEN_789;
  assign _GEN_791 = 11'h312 == _T_12323 ? mem_786 : _GEN_790;
  assign _GEN_792 = 11'h313 == _T_12323 ? mem_787 : _GEN_791;
  assign _GEN_793 = 11'h314 == _T_12323 ? mem_788 : _GEN_792;
  assign _GEN_794 = 11'h315 == _T_12323 ? mem_789 : _GEN_793;
  assign _GEN_795 = 11'h316 == _T_12323 ? mem_790 : _GEN_794;
  assign _GEN_796 = 11'h317 == _T_12323 ? mem_791 : _GEN_795;
  assign _GEN_797 = 11'h318 == _T_12323 ? mem_792 : _GEN_796;
  assign _GEN_798 = 11'h319 == _T_12323 ? mem_793 : _GEN_797;
  assign _GEN_799 = 11'h31a == _T_12323 ? mem_794 : _GEN_798;
  assign _GEN_800 = 11'h31b == _T_12323 ? mem_795 : _GEN_799;
  assign _GEN_801 = 11'h31c == _T_12323 ? mem_796 : _GEN_800;
  assign _GEN_802 = 11'h31d == _T_12323 ? mem_797 : _GEN_801;
  assign _GEN_803 = 11'h31e == _T_12323 ? mem_798 : _GEN_802;
  assign _GEN_804 = 11'h31f == _T_12323 ? mem_799 : _GEN_803;
  assign _GEN_805 = 11'h320 == _T_12323 ? mem_800 : _GEN_804;
  assign _GEN_806 = 11'h321 == _T_12323 ? mem_801 : _GEN_805;
  assign _GEN_807 = 11'h322 == _T_12323 ? mem_802 : _GEN_806;
  assign _GEN_808 = 11'h323 == _T_12323 ? mem_803 : _GEN_807;
  assign _GEN_809 = 11'h324 == _T_12323 ? mem_804 : _GEN_808;
  assign _GEN_810 = 11'h325 == _T_12323 ? mem_805 : _GEN_809;
  assign _GEN_811 = 11'h326 == _T_12323 ? mem_806 : _GEN_810;
  assign _GEN_812 = 11'h327 == _T_12323 ? mem_807 : _GEN_811;
  assign _GEN_813 = 11'h328 == _T_12323 ? mem_808 : _GEN_812;
  assign _GEN_814 = 11'h329 == _T_12323 ? mem_809 : _GEN_813;
  assign _GEN_815 = 11'h32a == _T_12323 ? mem_810 : _GEN_814;
  assign _GEN_816 = 11'h32b == _T_12323 ? mem_811 : _GEN_815;
  assign _GEN_817 = 11'h32c == _T_12323 ? mem_812 : _GEN_816;
  assign _GEN_818 = 11'h32d == _T_12323 ? mem_813 : _GEN_817;
  assign _GEN_819 = 11'h32e == _T_12323 ? mem_814 : _GEN_818;
  assign _GEN_820 = 11'h32f == _T_12323 ? mem_815 : _GEN_819;
  assign _GEN_821 = 11'h330 == _T_12323 ? mem_816 : _GEN_820;
  assign _GEN_822 = 11'h331 == _T_12323 ? mem_817 : _GEN_821;
  assign _GEN_823 = 11'h332 == _T_12323 ? mem_818 : _GEN_822;
  assign _GEN_824 = 11'h333 == _T_12323 ? mem_819 : _GEN_823;
  assign _GEN_825 = 11'h334 == _T_12323 ? mem_820 : _GEN_824;
  assign _GEN_826 = 11'h335 == _T_12323 ? mem_821 : _GEN_825;
  assign _GEN_827 = 11'h336 == _T_12323 ? mem_822 : _GEN_826;
  assign _GEN_828 = 11'h337 == _T_12323 ? mem_823 : _GEN_827;
  assign _GEN_829 = 11'h338 == _T_12323 ? mem_824 : _GEN_828;
  assign _GEN_830 = 11'h339 == _T_12323 ? mem_825 : _GEN_829;
  assign _GEN_831 = 11'h33a == _T_12323 ? mem_826 : _GEN_830;
  assign _GEN_832 = 11'h33b == _T_12323 ? mem_827 : _GEN_831;
  assign _GEN_833 = 11'h33c == _T_12323 ? mem_828 : _GEN_832;
  assign _GEN_834 = 11'h33d == _T_12323 ? mem_829 : _GEN_833;
  assign _GEN_835 = 11'h33e == _T_12323 ? mem_830 : _GEN_834;
  assign _GEN_836 = 11'h33f == _T_12323 ? mem_831 : _GEN_835;
  assign _GEN_837 = 11'h340 == _T_12323 ? mem_832 : _GEN_836;
  assign _GEN_838 = 11'h341 == _T_12323 ? mem_833 : _GEN_837;
  assign _GEN_839 = 11'h342 == _T_12323 ? mem_834 : _GEN_838;
  assign _GEN_840 = 11'h343 == _T_12323 ? mem_835 : _GEN_839;
  assign _GEN_841 = 11'h344 == _T_12323 ? mem_836 : _GEN_840;
  assign _GEN_842 = 11'h345 == _T_12323 ? mem_837 : _GEN_841;
  assign _GEN_843 = 11'h346 == _T_12323 ? mem_838 : _GEN_842;
  assign _GEN_844 = 11'h347 == _T_12323 ? mem_839 : _GEN_843;
  assign _GEN_845 = 11'h348 == _T_12323 ? mem_840 : _GEN_844;
  assign _GEN_846 = 11'h349 == _T_12323 ? mem_841 : _GEN_845;
  assign _GEN_847 = 11'h34a == _T_12323 ? mem_842 : _GEN_846;
  assign _GEN_848 = 11'h34b == _T_12323 ? mem_843 : _GEN_847;
  assign _GEN_849 = 11'h34c == _T_12323 ? mem_844 : _GEN_848;
  assign _GEN_850 = 11'h34d == _T_12323 ? mem_845 : _GEN_849;
  assign _GEN_851 = 11'h34e == _T_12323 ? mem_846 : _GEN_850;
  assign _GEN_852 = 11'h34f == _T_12323 ? mem_847 : _GEN_851;
  assign _GEN_853 = 11'h350 == _T_12323 ? mem_848 : _GEN_852;
  assign _GEN_854 = 11'h351 == _T_12323 ? mem_849 : _GEN_853;
  assign _GEN_855 = 11'h352 == _T_12323 ? mem_850 : _GEN_854;
  assign _GEN_856 = 11'h353 == _T_12323 ? mem_851 : _GEN_855;
  assign _GEN_857 = 11'h354 == _T_12323 ? mem_852 : _GEN_856;
  assign _GEN_858 = 11'h355 == _T_12323 ? mem_853 : _GEN_857;
  assign _GEN_859 = 11'h356 == _T_12323 ? mem_854 : _GEN_858;
  assign _GEN_860 = 11'h357 == _T_12323 ? mem_855 : _GEN_859;
  assign _GEN_861 = 11'h358 == _T_12323 ? mem_856 : _GEN_860;
  assign _GEN_862 = 11'h359 == _T_12323 ? mem_857 : _GEN_861;
  assign _GEN_863 = 11'h35a == _T_12323 ? mem_858 : _GEN_862;
  assign _GEN_864 = 11'h35b == _T_12323 ? mem_859 : _GEN_863;
  assign _GEN_865 = 11'h35c == _T_12323 ? mem_860 : _GEN_864;
  assign _GEN_866 = 11'h35d == _T_12323 ? mem_861 : _GEN_865;
  assign _GEN_867 = 11'h35e == _T_12323 ? mem_862 : _GEN_866;
  assign _GEN_868 = 11'h35f == _T_12323 ? mem_863 : _GEN_867;
  assign _GEN_869 = 11'h360 == _T_12323 ? mem_864 : _GEN_868;
  assign _GEN_870 = 11'h361 == _T_12323 ? mem_865 : _GEN_869;
  assign _GEN_871 = 11'h362 == _T_12323 ? mem_866 : _GEN_870;
  assign _GEN_872 = 11'h363 == _T_12323 ? mem_867 : _GEN_871;
  assign _GEN_873 = 11'h364 == _T_12323 ? mem_868 : _GEN_872;
  assign _GEN_874 = 11'h365 == _T_12323 ? mem_869 : _GEN_873;
  assign _GEN_875 = 11'h366 == _T_12323 ? mem_870 : _GEN_874;
  assign _GEN_876 = 11'h367 == _T_12323 ? mem_871 : _GEN_875;
  assign _GEN_877 = 11'h368 == _T_12323 ? mem_872 : _GEN_876;
  assign _GEN_878 = 11'h369 == _T_12323 ? mem_873 : _GEN_877;
  assign _GEN_879 = 11'h36a == _T_12323 ? mem_874 : _GEN_878;
  assign _GEN_880 = 11'h36b == _T_12323 ? mem_875 : _GEN_879;
  assign _GEN_881 = 11'h36c == _T_12323 ? mem_876 : _GEN_880;
  assign _GEN_882 = 11'h36d == _T_12323 ? mem_877 : _GEN_881;
  assign _GEN_883 = 11'h36e == _T_12323 ? mem_878 : _GEN_882;
  assign _GEN_884 = 11'h36f == _T_12323 ? mem_879 : _GEN_883;
  assign _GEN_885 = 11'h370 == _T_12323 ? mem_880 : _GEN_884;
  assign _GEN_886 = 11'h371 == _T_12323 ? mem_881 : _GEN_885;
  assign _GEN_887 = 11'h372 == _T_12323 ? mem_882 : _GEN_886;
  assign _GEN_888 = 11'h373 == _T_12323 ? mem_883 : _GEN_887;
  assign _GEN_889 = 11'h374 == _T_12323 ? mem_884 : _GEN_888;
  assign _GEN_890 = 11'h375 == _T_12323 ? mem_885 : _GEN_889;
  assign _GEN_891 = 11'h376 == _T_12323 ? mem_886 : _GEN_890;
  assign _GEN_892 = 11'h377 == _T_12323 ? mem_887 : _GEN_891;
  assign _GEN_893 = 11'h378 == _T_12323 ? mem_888 : _GEN_892;
  assign _GEN_894 = 11'h379 == _T_12323 ? mem_889 : _GEN_893;
  assign _GEN_895 = 11'h37a == _T_12323 ? mem_890 : _GEN_894;
  assign _GEN_896 = 11'h37b == _T_12323 ? mem_891 : _GEN_895;
  assign _GEN_897 = 11'h37c == _T_12323 ? mem_892 : _GEN_896;
  assign _GEN_898 = 11'h37d == _T_12323 ? mem_893 : _GEN_897;
  assign _GEN_899 = 11'h37e == _T_12323 ? mem_894 : _GEN_898;
  assign _GEN_900 = 11'h37f == _T_12323 ? mem_895 : _GEN_899;
  assign _GEN_901 = 11'h380 == _T_12323 ? mem_896 : _GEN_900;
  assign _GEN_902 = 11'h381 == _T_12323 ? mem_897 : _GEN_901;
  assign _GEN_903 = 11'h382 == _T_12323 ? mem_898 : _GEN_902;
  assign _GEN_904 = 11'h383 == _T_12323 ? mem_899 : _GEN_903;
  assign _GEN_905 = 11'h384 == _T_12323 ? mem_900 : _GEN_904;
  assign _GEN_906 = 11'h385 == _T_12323 ? mem_901 : _GEN_905;
  assign _GEN_907 = 11'h386 == _T_12323 ? mem_902 : _GEN_906;
  assign _GEN_908 = 11'h387 == _T_12323 ? mem_903 : _GEN_907;
  assign _GEN_909 = 11'h388 == _T_12323 ? mem_904 : _GEN_908;
  assign _GEN_910 = 11'h389 == _T_12323 ? mem_905 : _GEN_909;
  assign _GEN_911 = 11'h38a == _T_12323 ? mem_906 : _GEN_910;
  assign _GEN_912 = 11'h38b == _T_12323 ? mem_907 : _GEN_911;
  assign _GEN_913 = 11'h38c == _T_12323 ? mem_908 : _GEN_912;
  assign _GEN_914 = 11'h38d == _T_12323 ? mem_909 : _GEN_913;
  assign _GEN_915 = 11'h38e == _T_12323 ? mem_910 : _GEN_914;
  assign _GEN_916 = 11'h38f == _T_12323 ? mem_911 : _GEN_915;
  assign _GEN_917 = 11'h390 == _T_12323 ? mem_912 : _GEN_916;
  assign _GEN_918 = 11'h391 == _T_12323 ? mem_913 : _GEN_917;
  assign _GEN_919 = 11'h392 == _T_12323 ? mem_914 : _GEN_918;
  assign _GEN_920 = 11'h393 == _T_12323 ? mem_915 : _GEN_919;
  assign _GEN_921 = 11'h394 == _T_12323 ? mem_916 : _GEN_920;
  assign _GEN_922 = 11'h395 == _T_12323 ? mem_917 : _GEN_921;
  assign _GEN_923 = 11'h396 == _T_12323 ? mem_918 : _GEN_922;
  assign _GEN_924 = 11'h397 == _T_12323 ? mem_919 : _GEN_923;
  assign _GEN_925 = 11'h398 == _T_12323 ? mem_920 : _GEN_924;
  assign _GEN_926 = 11'h399 == _T_12323 ? mem_921 : _GEN_925;
  assign _GEN_927 = 11'h39a == _T_12323 ? mem_922 : _GEN_926;
  assign _GEN_928 = 11'h39b == _T_12323 ? mem_923 : _GEN_927;
  assign _GEN_929 = 11'h39c == _T_12323 ? mem_924 : _GEN_928;
  assign _GEN_930 = 11'h39d == _T_12323 ? mem_925 : _GEN_929;
  assign _GEN_931 = 11'h39e == _T_12323 ? mem_926 : _GEN_930;
  assign _GEN_932 = 11'h39f == _T_12323 ? mem_927 : _GEN_931;
  assign _GEN_933 = 11'h3a0 == _T_12323 ? mem_928 : _GEN_932;
  assign _GEN_934 = 11'h3a1 == _T_12323 ? mem_929 : _GEN_933;
  assign _GEN_935 = 11'h3a2 == _T_12323 ? mem_930 : _GEN_934;
  assign _GEN_936 = 11'h3a3 == _T_12323 ? mem_931 : _GEN_935;
  assign _GEN_937 = 11'h3a4 == _T_12323 ? mem_932 : _GEN_936;
  assign _GEN_938 = 11'h3a5 == _T_12323 ? mem_933 : _GEN_937;
  assign _GEN_939 = 11'h3a6 == _T_12323 ? mem_934 : _GEN_938;
  assign _GEN_940 = 11'h3a7 == _T_12323 ? mem_935 : _GEN_939;
  assign _GEN_941 = 11'h3a8 == _T_12323 ? mem_936 : _GEN_940;
  assign _GEN_942 = 11'h3a9 == _T_12323 ? mem_937 : _GEN_941;
  assign _GEN_943 = 11'h3aa == _T_12323 ? mem_938 : _GEN_942;
  assign _GEN_944 = 11'h3ab == _T_12323 ? mem_939 : _GEN_943;
  assign _GEN_945 = 11'h3ac == _T_12323 ? mem_940 : _GEN_944;
  assign _GEN_946 = 11'h3ad == _T_12323 ? mem_941 : _GEN_945;
  assign _GEN_947 = 11'h3ae == _T_12323 ? mem_942 : _GEN_946;
  assign _GEN_948 = 11'h3af == _T_12323 ? mem_943 : _GEN_947;
  assign _GEN_949 = 11'h3b0 == _T_12323 ? mem_944 : _GEN_948;
  assign _GEN_950 = 11'h3b1 == _T_12323 ? mem_945 : _GEN_949;
  assign _GEN_951 = 11'h3b2 == _T_12323 ? mem_946 : _GEN_950;
  assign _GEN_952 = 11'h3b3 == _T_12323 ? mem_947 : _GEN_951;
  assign _GEN_953 = 11'h3b4 == _T_12323 ? mem_948 : _GEN_952;
  assign _GEN_954 = 11'h3b5 == _T_12323 ? mem_949 : _GEN_953;
  assign _GEN_955 = 11'h3b6 == _T_12323 ? mem_950 : _GEN_954;
  assign _GEN_956 = 11'h3b7 == _T_12323 ? mem_951 : _GEN_955;
  assign _GEN_957 = 11'h3b8 == _T_12323 ? mem_952 : _GEN_956;
  assign _GEN_958 = 11'h3b9 == _T_12323 ? mem_953 : _GEN_957;
  assign _GEN_959 = 11'h3ba == _T_12323 ? mem_954 : _GEN_958;
  assign _GEN_960 = 11'h3bb == _T_12323 ? mem_955 : _GEN_959;
  assign _GEN_961 = 11'h3bc == _T_12323 ? mem_956 : _GEN_960;
  assign _GEN_962 = 11'h3bd == _T_12323 ? mem_957 : _GEN_961;
  assign _GEN_963 = 11'h3be == _T_12323 ? mem_958 : _GEN_962;
  assign _GEN_964 = 11'h3bf == _T_12323 ? mem_959 : _GEN_963;
  assign _GEN_965 = 11'h3c0 == _T_12323 ? mem_960 : _GEN_964;
  assign _GEN_966 = 11'h3c1 == _T_12323 ? mem_961 : _GEN_965;
  assign _GEN_967 = 11'h3c2 == _T_12323 ? mem_962 : _GEN_966;
  assign _GEN_968 = 11'h3c3 == _T_12323 ? mem_963 : _GEN_967;
  assign _GEN_969 = 11'h3c4 == _T_12323 ? mem_964 : _GEN_968;
  assign _GEN_970 = 11'h3c5 == _T_12323 ? mem_965 : _GEN_969;
  assign _GEN_971 = 11'h3c6 == _T_12323 ? mem_966 : _GEN_970;
  assign _GEN_972 = 11'h3c7 == _T_12323 ? mem_967 : _GEN_971;
  assign _GEN_973 = 11'h3c8 == _T_12323 ? mem_968 : _GEN_972;
  assign _GEN_974 = 11'h3c9 == _T_12323 ? mem_969 : _GEN_973;
  assign _GEN_975 = 11'h3ca == _T_12323 ? mem_970 : _GEN_974;
  assign _GEN_976 = 11'h3cb == _T_12323 ? mem_971 : _GEN_975;
  assign _GEN_977 = 11'h3cc == _T_12323 ? mem_972 : _GEN_976;
  assign _GEN_978 = 11'h3cd == _T_12323 ? mem_973 : _GEN_977;
  assign _GEN_979 = 11'h3ce == _T_12323 ? mem_974 : _GEN_978;
  assign _GEN_980 = 11'h3cf == _T_12323 ? mem_975 : _GEN_979;
  assign _GEN_981 = 11'h3d0 == _T_12323 ? mem_976 : _GEN_980;
  assign _GEN_982 = 11'h3d1 == _T_12323 ? mem_977 : _GEN_981;
  assign _GEN_983 = 11'h3d2 == _T_12323 ? mem_978 : _GEN_982;
  assign _GEN_984 = 11'h3d3 == _T_12323 ? mem_979 : _GEN_983;
  assign _GEN_985 = 11'h3d4 == _T_12323 ? mem_980 : _GEN_984;
  assign _GEN_986 = 11'h3d5 == _T_12323 ? mem_981 : _GEN_985;
  assign _GEN_987 = 11'h3d6 == _T_12323 ? mem_982 : _GEN_986;
  assign _GEN_988 = 11'h3d7 == _T_12323 ? mem_983 : _GEN_987;
  assign _GEN_989 = 11'h3d8 == _T_12323 ? mem_984 : _GEN_988;
  assign _GEN_990 = 11'h3d9 == _T_12323 ? mem_985 : _GEN_989;
  assign _GEN_991 = 11'h3da == _T_12323 ? mem_986 : _GEN_990;
  assign _GEN_992 = 11'h3db == _T_12323 ? mem_987 : _GEN_991;
  assign _GEN_993 = 11'h3dc == _T_12323 ? mem_988 : _GEN_992;
  assign _GEN_994 = 11'h3dd == _T_12323 ? mem_989 : _GEN_993;
  assign _GEN_995 = 11'h3de == _T_12323 ? mem_990 : _GEN_994;
  assign _GEN_996 = 11'h3df == _T_12323 ? mem_991 : _GEN_995;
  assign _GEN_997 = 11'h3e0 == _T_12323 ? mem_992 : _GEN_996;
  assign _GEN_998 = 11'h3e1 == _T_12323 ? mem_993 : _GEN_997;
  assign _GEN_999 = 11'h3e2 == _T_12323 ? mem_994 : _GEN_998;
  assign _GEN_1000 = 11'h3e3 == _T_12323 ? mem_995 : _GEN_999;
  assign _GEN_1001 = 11'h3e4 == _T_12323 ? mem_996 : _GEN_1000;
  assign _GEN_1002 = 11'h3e5 == _T_12323 ? mem_997 : _GEN_1001;
  assign _GEN_1003 = 11'h3e6 == _T_12323 ? mem_998 : _GEN_1002;
  assign _GEN_1004 = 11'h3e7 == _T_12323 ? mem_999 : _GEN_1003;
  assign _GEN_1005 = 11'h3e8 == _T_12323 ? mem_1000 : _GEN_1004;
  assign _GEN_1006 = 11'h3e9 == _T_12323 ? mem_1001 : _GEN_1005;
  assign _GEN_1007 = 11'h3ea == _T_12323 ? mem_1002 : _GEN_1006;
  assign _GEN_1008 = 11'h3eb == _T_12323 ? mem_1003 : _GEN_1007;
  assign _GEN_1009 = 11'h3ec == _T_12323 ? mem_1004 : _GEN_1008;
  assign _GEN_1010 = 11'h3ed == _T_12323 ? mem_1005 : _GEN_1009;
  assign _GEN_1011 = 11'h3ee == _T_12323 ? mem_1006 : _GEN_1010;
  assign _GEN_1012 = 11'h3ef == _T_12323 ? mem_1007 : _GEN_1011;
  assign _GEN_1013 = 11'h3f0 == _T_12323 ? mem_1008 : _GEN_1012;
  assign _GEN_1014 = 11'h3f1 == _T_12323 ? mem_1009 : _GEN_1013;
  assign _GEN_1015 = 11'h3f2 == _T_12323 ? mem_1010 : _GEN_1014;
  assign _GEN_1016 = 11'h3f3 == _T_12323 ? mem_1011 : _GEN_1015;
  assign _GEN_1017 = 11'h3f4 == _T_12323 ? mem_1012 : _GEN_1016;
  assign _GEN_1018 = 11'h3f5 == _T_12323 ? mem_1013 : _GEN_1017;
  assign _GEN_1019 = 11'h3f6 == _T_12323 ? mem_1014 : _GEN_1018;
  assign _GEN_1020 = 11'h3f7 == _T_12323 ? mem_1015 : _GEN_1019;
  assign _GEN_1021 = 11'h3f8 == _T_12323 ? mem_1016 : _GEN_1020;
  assign _GEN_1022 = 11'h3f9 == _T_12323 ? mem_1017 : _GEN_1021;
  assign _GEN_1023 = 11'h3fa == _T_12323 ? mem_1018 : _GEN_1022;
  assign _GEN_1024 = 11'h3fb == _T_12323 ? mem_1019 : _GEN_1023;
  assign _GEN_1025 = 11'h3fc == _T_12323 ? mem_1020 : _GEN_1024;
  assign _GEN_1026 = 11'h3fd == _T_12323 ? mem_1021 : _GEN_1025;
  assign _GEN_1027 = 11'h3fe == _T_12323 ? mem_1022 : _GEN_1026;
  assign _GEN_1028 = 11'h3ff == _T_12323 ? mem_1023 : _GEN_1027;
  assign _GEN_1029 = 11'h400 == _T_12323 ? mem_1024 : _GEN_1028;
  assign _GEN_1030 = 11'h401 == _T_12323 ? mem_1025 : _GEN_1029;
  assign _GEN_1031 = 11'h402 == _T_12323 ? mem_1026 : _GEN_1030;
  assign _GEN_1032 = 11'h403 == _T_12323 ? mem_1027 : _GEN_1031;
  assign _GEN_1033 = 11'h404 == _T_12323 ? mem_1028 : _GEN_1032;
  assign _GEN_1034 = 11'h405 == _T_12323 ? mem_1029 : _GEN_1033;
  assign _GEN_1035 = 11'h406 == _T_12323 ? mem_1030 : _GEN_1034;
  assign _GEN_1036 = 11'h407 == _T_12323 ? mem_1031 : _GEN_1035;
  assign _GEN_1037 = 11'h408 == _T_12323 ? mem_1032 : _GEN_1036;
  assign _GEN_1038 = 11'h409 == _T_12323 ? mem_1033 : _GEN_1037;
  assign _GEN_1039 = 11'h40a == _T_12323 ? mem_1034 : _GEN_1038;
  assign _GEN_1040 = 11'h40b == _T_12323 ? mem_1035 : _GEN_1039;
  assign _GEN_1041 = 11'h40c == _T_12323 ? mem_1036 : _GEN_1040;
  assign _GEN_1042 = 11'h40d == _T_12323 ? mem_1037 : _GEN_1041;
  assign _GEN_1043 = 11'h40e == _T_12323 ? mem_1038 : _GEN_1042;
  assign _GEN_1044 = 11'h40f == _T_12323 ? mem_1039 : _GEN_1043;
  assign _GEN_1045 = 11'h410 == _T_12323 ? mem_1040 : _GEN_1044;
  assign _GEN_1046 = 11'h411 == _T_12323 ? mem_1041 : _GEN_1045;
  assign _GEN_1047 = 11'h412 == _T_12323 ? mem_1042 : _GEN_1046;
  assign _GEN_1048 = 11'h413 == _T_12323 ? mem_1043 : _GEN_1047;
  assign _GEN_1049 = 11'h414 == _T_12323 ? mem_1044 : _GEN_1048;
  assign _GEN_1050 = 11'h415 == _T_12323 ? mem_1045 : _GEN_1049;
  assign _GEN_1051 = 11'h416 == _T_12323 ? mem_1046 : _GEN_1050;
  assign _GEN_1052 = 11'h417 == _T_12323 ? mem_1047 : _GEN_1051;
  assign _GEN_1053 = 11'h418 == _T_12323 ? mem_1048 : _GEN_1052;
  assign _GEN_1054 = 11'h419 == _T_12323 ? mem_1049 : _GEN_1053;
  assign _GEN_1055 = 11'h41a == _T_12323 ? mem_1050 : _GEN_1054;
  assign _GEN_1056 = 11'h41b == _T_12323 ? mem_1051 : _GEN_1055;
  assign _GEN_1057 = 11'h41c == _T_12323 ? mem_1052 : _GEN_1056;
  assign _GEN_1058 = 11'h41d == _T_12323 ? mem_1053 : _GEN_1057;
  assign _GEN_1059 = 11'h41e == _T_12323 ? mem_1054 : _GEN_1058;
  assign _GEN_1060 = 11'h41f == _T_12323 ? mem_1055 : _GEN_1059;
  assign _GEN_1061 = 11'h420 == _T_12323 ? mem_1056 : _GEN_1060;
  assign _GEN_1062 = 11'h421 == _T_12323 ? mem_1057 : _GEN_1061;
  assign _GEN_1063 = 11'h422 == _T_12323 ? mem_1058 : _GEN_1062;
  assign _GEN_1064 = 11'h423 == _T_12323 ? mem_1059 : _GEN_1063;
  assign _GEN_1065 = 11'h424 == _T_12323 ? mem_1060 : _GEN_1064;
  assign _GEN_1066 = 11'h425 == _T_12323 ? mem_1061 : _GEN_1065;
  assign _GEN_1067 = 11'h426 == _T_12323 ? mem_1062 : _GEN_1066;
  assign _GEN_1068 = 11'h427 == _T_12323 ? mem_1063 : _GEN_1067;
  assign _GEN_1069 = 11'h428 == _T_12323 ? mem_1064 : _GEN_1068;
  assign _GEN_1070 = 11'h429 == _T_12323 ? mem_1065 : _GEN_1069;
  assign _GEN_1071 = 11'h42a == _T_12323 ? mem_1066 : _GEN_1070;
  assign _GEN_1072 = 11'h42b == _T_12323 ? mem_1067 : _GEN_1071;
  assign _GEN_1073 = 11'h42c == _T_12323 ? mem_1068 : _GEN_1072;
  assign _GEN_1074 = 11'h42d == _T_12323 ? mem_1069 : _GEN_1073;
  assign _GEN_1075 = 11'h42e == _T_12323 ? mem_1070 : _GEN_1074;
  assign _GEN_1076 = 11'h42f == _T_12323 ? mem_1071 : _GEN_1075;
  assign _GEN_1077 = 11'h430 == _T_12323 ? mem_1072 : _GEN_1076;
  assign _GEN_1078 = 11'h431 == _T_12323 ? mem_1073 : _GEN_1077;
  assign _GEN_1079 = 11'h432 == _T_12323 ? mem_1074 : _GEN_1078;
  assign _GEN_1080 = 11'h433 == _T_12323 ? mem_1075 : _GEN_1079;
  assign _GEN_1081 = 11'h434 == _T_12323 ? mem_1076 : _GEN_1080;
  assign _GEN_1082 = 11'h435 == _T_12323 ? mem_1077 : _GEN_1081;
  assign _GEN_1083 = 11'h436 == _T_12323 ? mem_1078 : _GEN_1082;
  assign _GEN_1084 = 11'h437 == _T_12323 ? mem_1079 : _GEN_1083;
  assign _GEN_1085 = 11'h438 == _T_12323 ? mem_1080 : _GEN_1084;
  assign _GEN_1086 = 11'h439 == _T_12323 ? mem_1081 : _GEN_1085;
  assign _GEN_1087 = 11'h43a == _T_12323 ? mem_1082 : _GEN_1086;
  assign _GEN_1088 = 11'h43b == _T_12323 ? mem_1083 : _GEN_1087;
  assign _GEN_1089 = 11'h43c == _T_12323 ? mem_1084 : _GEN_1088;
  assign _GEN_1090 = 11'h43d == _T_12323 ? mem_1085 : _GEN_1089;
  assign _GEN_1091 = 11'h43e == _T_12323 ? mem_1086 : _GEN_1090;
  assign _GEN_1092 = 11'h43f == _T_12323 ? mem_1087 : _GEN_1091;
  assign _GEN_1093 = 11'h440 == _T_12323 ? mem_1088 : _GEN_1092;
  assign _GEN_1094 = 11'h441 == _T_12323 ? mem_1089 : _GEN_1093;
  assign _GEN_1095 = 11'h442 == _T_12323 ? mem_1090 : _GEN_1094;
  assign _GEN_1096 = 11'h443 == _T_12323 ? mem_1091 : _GEN_1095;
  assign _GEN_1097 = 11'h444 == _T_12323 ? mem_1092 : _GEN_1096;
  assign _GEN_1098 = 11'h445 == _T_12323 ? mem_1093 : _GEN_1097;
  assign _GEN_1099 = 11'h446 == _T_12323 ? mem_1094 : _GEN_1098;
  assign _GEN_1100 = 11'h447 == _T_12323 ? mem_1095 : _GEN_1099;
  assign _GEN_1101 = 11'h448 == _T_12323 ? mem_1096 : _GEN_1100;
  assign _GEN_1102 = 11'h449 == _T_12323 ? mem_1097 : _GEN_1101;
  assign _GEN_1103 = 11'h44a == _T_12323 ? mem_1098 : _GEN_1102;
  assign _GEN_1104 = 11'h44b == _T_12323 ? mem_1099 : _GEN_1103;
  assign _GEN_1105 = 11'h44c == _T_12323 ? mem_1100 : _GEN_1104;
  assign _GEN_1106 = 11'h44d == _T_12323 ? mem_1101 : _GEN_1105;
  assign _GEN_1107 = 11'h44e == _T_12323 ? mem_1102 : _GEN_1106;
  assign _GEN_1108 = 11'h44f == _T_12323 ? mem_1103 : _GEN_1107;
  assign _GEN_1109 = 11'h450 == _T_12323 ? mem_1104 : _GEN_1108;
  assign _GEN_1110 = 11'h451 == _T_12323 ? mem_1105 : _GEN_1109;
  assign _GEN_1111 = 11'h452 == _T_12323 ? mem_1106 : _GEN_1110;
  assign _GEN_1112 = 11'h453 == _T_12323 ? mem_1107 : _GEN_1111;
  assign _GEN_1113 = 11'h454 == _T_12323 ? mem_1108 : _GEN_1112;
  assign _GEN_1114 = 11'h455 == _T_12323 ? mem_1109 : _GEN_1113;
  assign _GEN_1115 = 11'h456 == _T_12323 ? mem_1110 : _GEN_1114;
  assign _GEN_1116 = 11'h457 == _T_12323 ? mem_1111 : _GEN_1115;
  assign _GEN_1117 = 11'h458 == _T_12323 ? mem_1112 : _GEN_1116;
  assign _GEN_1118 = 11'h459 == _T_12323 ? mem_1113 : _GEN_1117;
  assign _GEN_1119 = 11'h45a == _T_12323 ? mem_1114 : _GEN_1118;
  assign _GEN_1120 = 11'h45b == _T_12323 ? mem_1115 : _GEN_1119;
  assign _GEN_1121 = 11'h45c == _T_12323 ? mem_1116 : _GEN_1120;
  assign _GEN_1122 = 11'h45d == _T_12323 ? mem_1117 : _GEN_1121;
  assign _GEN_1123 = 11'h45e == _T_12323 ? mem_1118 : _GEN_1122;
  assign _GEN_1124 = 11'h45f == _T_12323 ? mem_1119 : _GEN_1123;
  assign _GEN_1125 = 11'h460 == _T_12323 ? mem_1120 : _GEN_1124;
  assign _GEN_1126 = 11'h461 == _T_12323 ? mem_1121 : _GEN_1125;
  assign _GEN_1127 = 11'h462 == _T_12323 ? mem_1122 : _GEN_1126;
  assign _GEN_1128 = 11'h463 == _T_12323 ? mem_1123 : _GEN_1127;
  assign _GEN_1129 = 11'h464 == _T_12323 ? mem_1124 : _GEN_1128;
  assign _GEN_1130 = 11'h465 == _T_12323 ? mem_1125 : _GEN_1129;
  assign _GEN_1131 = 11'h466 == _T_12323 ? mem_1126 : _GEN_1130;
  assign _GEN_1132 = 11'h467 == _T_12323 ? mem_1127 : _GEN_1131;
  assign _GEN_1133 = 11'h468 == _T_12323 ? mem_1128 : _GEN_1132;
  assign _GEN_1134 = 11'h469 == _T_12323 ? mem_1129 : _GEN_1133;
  assign _GEN_1135 = 11'h46a == _T_12323 ? mem_1130 : _GEN_1134;
  assign _GEN_1136 = 11'h46b == _T_12323 ? mem_1131 : _GEN_1135;
  assign _GEN_1137 = 11'h46c == _T_12323 ? mem_1132 : _GEN_1136;
  assign _GEN_1138 = 11'h46d == _T_12323 ? mem_1133 : _GEN_1137;
  assign _GEN_1139 = 11'h46e == _T_12323 ? mem_1134 : _GEN_1138;
  assign _GEN_1140 = 11'h46f == _T_12323 ? mem_1135 : _GEN_1139;
  assign _GEN_1141 = 11'h470 == _T_12323 ? mem_1136 : _GEN_1140;
  assign _GEN_1142 = 11'h471 == _T_12323 ? mem_1137 : _GEN_1141;
  assign _GEN_1143 = 11'h472 == _T_12323 ? mem_1138 : _GEN_1142;
  assign _GEN_1144 = 11'h473 == _T_12323 ? mem_1139 : _GEN_1143;
  assign _GEN_1145 = 11'h474 == _T_12323 ? mem_1140 : _GEN_1144;
  assign _GEN_1146 = 11'h475 == _T_12323 ? mem_1141 : _GEN_1145;
  assign _GEN_1147 = 11'h476 == _T_12323 ? mem_1142 : _GEN_1146;
  assign _GEN_1148 = 11'h477 == _T_12323 ? mem_1143 : _GEN_1147;
  assign _GEN_1149 = 11'h478 == _T_12323 ? mem_1144 : _GEN_1148;
  assign _GEN_1150 = 11'h479 == _T_12323 ? mem_1145 : _GEN_1149;
  assign _GEN_1151 = 11'h47a == _T_12323 ? mem_1146 : _GEN_1150;
  assign _GEN_1152 = 11'h47b == _T_12323 ? mem_1147 : _GEN_1151;
  assign _GEN_1153 = 11'h47c == _T_12323 ? mem_1148 : _GEN_1152;
  assign _GEN_1154 = 11'h47d == _T_12323 ? mem_1149 : _GEN_1153;
  assign _GEN_1155 = 11'h47e == _T_12323 ? mem_1150 : _GEN_1154;
  assign _GEN_1156 = 11'h47f == _T_12323 ? mem_1151 : _GEN_1155;
  assign _GEN_1157 = 11'h480 == _T_12323 ? mem_1152 : _GEN_1156;
  assign _GEN_1158 = 11'h481 == _T_12323 ? mem_1153 : _GEN_1157;
  assign _GEN_1159 = 11'h482 == _T_12323 ? mem_1154 : _GEN_1158;
  assign _GEN_1160 = 11'h483 == _T_12323 ? mem_1155 : _GEN_1159;
  assign _GEN_1161 = 11'h484 == _T_12323 ? mem_1156 : _GEN_1160;
  assign _GEN_1162 = 11'h485 == _T_12323 ? mem_1157 : _GEN_1161;
  assign _GEN_1163 = 11'h486 == _T_12323 ? mem_1158 : _GEN_1162;
  assign _GEN_1164 = 11'h487 == _T_12323 ? mem_1159 : _GEN_1163;
  assign _GEN_1165 = 11'h488 == _T_12323 ? mem_1160 : _GEN_1164;
  assign _GEN_1166 = 11'h489 == _T_12323 ? mem_1161 : _GEN_1165;
  assign _GEN_1167 = 11'h48a == _T_12323 ? mem_1162 : _GEN_1166;
  assign _GEN_1168 = 11'h48b == _T_12323 ? mem_1163 : _GEN_1167;
  assign _GEN_1169 = 11'h48c == _T_12323 ? mem_1164 : _GEN_1168;
  assign _GEN_1170 = 11'h48d == _T_12323 ? mem_1165 : _GEN_1169;
  assign _GEN_1171 = 11'h48e == _T_12323 ? mem_1166 : _GEN_1170;
  assign _GEN_1172 = 11'h48f == _T_12323 ? mem_1167 : _GEN_1171;
  assign _GEN_1173 = 11'h490 == _T_12323 ? mem_1168 : _GEN_1172;
  assign _GEN_1174 = 11'h491 == _T_12323 ? mem_1169 : _GEN_1173;
  assign _GEN_1175 = 11'h492 == _T_12323 ? mem_1170 : _GEN_1174;
  assign _GEN_1176 = 11'h493 == _T_12323 ? mem_1171 : _GEN_1175;
  assign _GEN_1177 = 11'h494 == _T_12323 ? mem_1172 : _GEN_1176;
  assign _GEN_1178 = 11'h495 == _T_12323 ? mem_1173 : _GEN_1177;
  assign _GEN_1179 = 11'h496 == _T_12323 ? mem_1174 : _GEN_1178;
  assign _GEN_1180 = 11'h497 == _T_12323 ? mem_1175 : _GEN_1179;
  assign _GEN_1181 = 11'h498 == _T_12323 ? mem_1176 : _GEN_1180;
  assign _GEN_1182 = 11'h499 == _T_12323 ? mem_1177 : _GEN_1181;
  assign _GEN_1183 = 11'h49a == _T_12323 ? mem_1178 : _GEN_1182;
  assign _GEN_1184 = 11'h49b == _T_12323 ? mem_1179 : _GEN_1183;
  assign _GEN_1185 = 11'h49c == _T_12323 ? mem_1180 : _GEN_1184;
  assign _GEN_1186 = 11'h49d == _T_12323 ? mem_1181 : _GEN_1185;
  assign _GEN_1187 = 11'h49e == _T_12323 ? mem_1182 : _GEN_1186;
  assign _GEN_1188 = 11'h49f == _T_12323 ? mem_1183 : _GEN_1187;
  assign _GEN_1189 = 11'h4a0 == _T_12323 ? mem_1184 : _GEN_1188;
  assign _GEN_1190 = 11'h4a1 == _T_12323 ? mem_1185 : _GEN_1189;
  assign _GEN_1191 = 11'h4a2 == _T_12323 ? mem_1186 : _GEN_1190;
  assign _GEN_1192 = 11'h4a3 == _T_12323 ? mem_1187 : _GEN_1191;
  assign _GEN_1193 = 11'h4a4 == _T_12323 ? mem_1188 : _GEN_1192;
  assign _GEN_1194 = 11'h4a5 == _T_12323 ? mem_1189 : _GEN_1193;
  assign _GEN_1195 = 11'h4a6 == _T_12323 ? mem_1190 : _GEN_1194;
  assign _GEN_1196 = 11'h4a7 == _T_12323 ? mem_1191 : _GEN_1195;
  assign _GEN_1197 = 11'h4a8 == _T_12323 ? mem_1192 : _GEN_1196;
  assign _GEN_1198 = 11'h4a9 == _T_12323 ? mem_1193 : _GEN_1197;
  assign _GEN_1199 = 11'h4aa == _T_12323 ? mem_1194 : _GEN_1198;
  assign _GEN_1200 = 11'h4ab == _T_12323 ? mem_1195 : _GEN_1199;
  assign _GEN_1201 = 11'h4ac == _T_12323 ? mem_1196 : _GEN_1200;
  assign _GEN_1202 = 11'h4ad == _T_12323 ? mem_1197 : _GEN_1201;
  assign _GEN_1203 = 11'h4ae == _T_12323 ? mem_1198 : _GEN_1202;
  assign _GEN_1204 = 11'h4af == _T_12323 ? mem_1199 : _GEN_1203;
  assign _GEN_1205 = 11'h4b0 == _T_12323 ? mem_1200 : _GEN_1204;
  assign _GEN_1206 = 11'h4b1 == _T_12323 ? mem_1201 : _GEN_1205;
  assign _GEN_1207 = 11'h4b2 == _T_12323 ? mem_1202 : _GEN_1206;
  assign _GEN_1208 = 11'h4b3 == _T_12323 ? mem_1203 : _GEN_1207;
  assign _GEN_1209 = 11'h4b4 == _T_12323 ? mem_1204 : _GEN_1208;
  assign _GEN_1210 = 11'h4b5 == _T_12323 ? mem_1205 : _GEN_1209;
  assign _GEN_1211 = 11'h4b6 == _T_12323 ? mem_1206 : _GEN_1210;
  assign _GEN_1212 = 11'h4b7 == _T_12323 ? mem_1207 : _GEN_1211;
  assign _GEN_1213 = 11'h4b8 == _T_12323 ? mem_1208 : _GEN_1212;
  assign _GEN_1214 = 11'h4b9 == _T_12323 ? mem_1209 : _GEN_1213;
  assign _GEN_1215 = 11'h4ba == _T_12323 ? mem_1210 : _GEN_1214;
  assign _GEN_1216 = 11'h4bb == _T_12323 ? mem_1211 : _GEN_1215;
  assign _GEN_1217 = 11'h4bc == _T_12323 ? mem_1212 : _GEN_1216;
  assign _GEN_1218 = 11'h4bd == _T_12323 ? mem_1213 : _GEN_1217;
  assign _GEN_1219 = 11'h4be == _T_12323 ? mem_1214 : _GEN_1218;
  assign _GEN_1220 = 11'h4bf == _T_12323 ? mem_1215 : _GEN_1219;
  assign _GEN_1221 = 11'h4c0 == _T_12323 ? mem_1216 : _GEN_1220;
  assign _GEN_1222 = 11'h4c1 == _T_12323 ? mem_1217 : _GEN_1221;
  assign _GEN_1223 = 11'h4c2 == _T_12323 ? mem_1218 : _GEN_1222;
  assign _GEN_1224 = 11'h4c3 == _T_12323 ? mem_1219 : _GEN_1223;
  assign _GEN_1225 = 11'h4c4 == _T_12323 ? mem_1220 : _GEN_1224;
  assign _GEN_1226 = 11'h4c5 == _T_12323 ? mem_1221 : _GEN_1225;
  assign _GEN_1227 = 11'h4c6 == _T_12323 ? mem_1222 : _GEN_1226;
  assign _GEN_1228 = 11'h4c7 == _T_12323 ? mem_1223 : _GEN_1227;
  assign _GEN_1229 = 11'h4c8 == _T_12323 ? mem_1224 : _GEN_1228;
  assign _GEN_1230 = 11'h4c9 == _T_12323 ? mem_1225 : _GEN_1229;
  assign _GEN_1231 = 11'h4ca == _T_12323 ? mem_1226 : _GEN_1230;
  assign _GEN_1232 = 11'h4cb == _T_12323 ? mem_1227 : _GEN_1231;
  assign _GEN_1233 = 11'h4cc == _T_12323 ? mem_1228 : _GEN_1232;
  assign _GEN_1234 = 11'h4cd == _T_12323 ? mem_1229 : _GEN_1233;
  assign _GEN_1235 = 11'h4ce == _T_12323 ? mem_1230 : _GEN_1234;
  assign _GEN_1236 = 11'h4cf == _T_12323 ? mem_1231 : _GEN_1235;
  assign _GEN_1237 = 11'h4d0 == _T_12323 ? mem_1232 : _GEN_1236;
  assign _GEN_1238 = 11'h4d1 == _T_12323 ? mem_1233 : _GEN_1237;
  assign _GEN_1239 = 11'h4d2 == _T_12323 ? mem_1234 : _GEN_1238;
  assign _GEN_1240 = 11'h4d3 == _T_12323 ? mem_1235 : _GEN_1239;
  assign _GEN_1241 = 11'h4d4 == _T_12323 ? mem_1236 : _GEN_1240;
  assign _GEN_1242 = 11'h4d5 == _T_12323 ? mem_1237 : _GEN_1241;
  assign _GEN_1243 = 11'h4d6 == _T_12323 ? mem_1238 : _GEN_1242;
  assign _GEN_1244 = 11'h4d7 == _T_12323 ? mem_1239 : _GEN_1243;
  assign _GEN_1245 = 11'h4d8 == _T_12323 ? mem_1240 : _GEN_1244;
  assign _GEN_1246 = 11'h4d9 == _T_12323 ? mem_1241 : _GEN_1245;
  assign _GEN_1247 = 11'h4da == _T_12323 ? mem_1242 : _GEN_1246;
  assign _GEN_1248 = 11'h4db == _T_12323 ? mem_1243 : _GEN_1247;
  assign _GEN_1249 = 11'h4dc == _T_12323 ? mem_1244 : _GEN_1248;
  assign _GEN_1250 = 11'h4dd == _T_12323 ? mem_1245 : _GEN_1249;
  assign _GEN_1251 = 11'h4de == _T_12323 ? mem_1246 : _GEN_1250;
  assign _GEN_1252 = 11'h4df == _T_12323 ? mem_1247 : _GEN_1251;
  assign _GEN_1253 = 11'h4e0 == _T_12323 ? mem_1248 : _GEN_1252;
  assign _GEN_1254 = 11'h4e1 == _T_12323 ? mem_1249 : _GEN_1253;
  assign _GEN_1255 = 11'h4e2 == _T_12323 ? mem_1250 : _GEN_1254;
  assign _GEN_1256 = 11'h4e3 == _T_12323 ? mem_1251 : _GEN_1255;
  assign _GEN_1257 = 11'h4e4 == _T_12323 ? mem_1252 : _GEN_1256;
  assign _GEN_1258 = 11'h4e5 == _T_12323 ? mem_1253 : _GEN_1257;
  assign _GEN_1259 = 11'h4e6 == _T_12323 ? mem_1254 : _GEN_1258;
  assign _GEN_1260 = 11'h4e7 == _T_12323 ? mem_1255 : _GEN_1259;
  assign _GEN_1261 = 11'h4e8 == _T_12323 ? mem_1256 : _GEN_1260;
  assign _GEN_1262 = 11'h4e9 == _T_12323 ? mem_1257 : _GEN_1261;
  assign _GEN_1263 = 11'h4ea == _T_12323 ? mem_1258 : _GEN_1262;
  assign _GEN_1264 = 11'h4eb == _T_12323 ? mem_1259 : _GEN_1263;
  assign _GEN_1265 = 11'h4ec == _T_12323 ? mem_1260 : _GEN_1264;
  assign _GEN_1266 = 11'h4ed == _T_12323 ? mem_1261 : _GEN_1265;
  assign _GEN_1267 = 11'h4ee == _T_12323 ? mem_1262 : _GEN_1266;
  assign _GEN_1268 = 11'h4ef == _T_12323 ? mem_1263 : _GEN_1267;
  assign _GEN_1269 = 11'h4f0 == _T_12323 ? mem_1264 : _GEN_1268;
  assign _GEN_1270 = 11'h4f1 == _T_12323 ? mem_1265 : _GEN_1269;
  assign _GEN_1271 = 11'h4f2 == _T_12323 ? mem_1266 : _GEN_1270;
  assign _GEN_1272 = 11'h4f3 == _T_12323 ? mem_1267 : _GEN_1271;
  assign _GEN_1273 = 11'h4f4 == _T_12323 ? mem_1268 : _GEN_1272;
  assign _GEN_1274 = 11'h4f5 == _T_12323 ? mem_1269 : _GEN_1273;
  assign _GEN_1275 = 11'h4f6 == _T_12323 ? mem_1270 : _GEN_1274;
  assign _GEN_1276 = 11'h4f7 == _T_12323 ? mem_1271 : _GEN_1275;
  assign _GEN_1277 = 11'h4f8 == _T_12323 ? mem_1272 : _GEN_1276;
  assign _GEN_1278 = 11'h4f9 == _T_12323 ? mem_1273 : _GEN_1277;
  assign _GEN_1279 = 11'h4fa == _T_12323 ? mem_1274 : _GEN_1278;
  assign _GEN_1280 = 11'h4fb == _T_12323 ? mem_1275 : _GEN_1279;
  assign _GEN_1281 = 11'h4fc == _T_12323 ? mem_1276 : _GEN_1280;
  assign _GEN_1282 = 11'h4fd == _T_12323 ? mem_1277 : _GEN_1281;
  assign _GEN_1283 = 11'h4fe == _T_12323 ? mem_1278 : _GEN_1282;
  assign _GEN_1284 = 11'h4ff == _T_12323 ? mem_1279 : _GEN_1283;
  assign _GEN_1285 = 11'h500 == _T_12323 ? mem_1280 : _GEN_1284;
  assign _GEN_1286 = 11'h501 == _T_12323 ? mem_1281 : _GEN_1285;
  assign _GEN_1287 = 11'h502 == _T_12323 ? mem_1282 : _GEN_1286;
  assign _GEN_1288 = 11'h503 == _T_12323 ? mem_1283 : _GEN_1287;
  assign _GEN_1289 = 11'h504 == _T_12323 ? mem_1284 : _GEN_1288;
  assign _GEN_1290 = 11'h505 == _T_12323 ? mem_1285 : _GEN_1289;
  assign _GEN_1291 = 11'h506 == _T_12323 ? mem_1286 : _GEN_1290;
  assign _GEN_1292 = 11'h507 == _T_12323 ? mem_1287 : _GEN_1291;
  assign _GEN_1293 = 11'h508 == _T_12323 ? mem_1288 : _GEN_1292;
  assign _GEN_1294 = 11'h509 == _T_12323 ? mem_1289 : _GEN_1293;
  assign _GEN_1295 = 11'h50a == _T_12323 ? mem_1290 : _GEN_1294;
  assign _GEN_1296 = 11'h50b == _T_12323 ? mem_1291 : _GEN_1295;
  assign _GEN_1297 = 11'h50c == _T_12323 ? mem_1292 : _GEN_1296;
  assign _GEN_1298 = 11'h50d == _T_12323 ? mem_1293 : _GEN_1297;
  assign _GEN_1299 = 11'h50e == _T_12323 ? mem_1294 : _GEN_1298;
  assign _GEN_1300 = 11'h50f == _T_12323 ? mem_1295 : _GEN_1299;
  assign _GEN_1301 = 11'h510 == _T_12323 ? mem_1296 : _GEN_1300;
  assign _GEN_1302 = 11'h511 == _T_12323 ? mem_1297 : _GEN_1301;
  assign _GEN_1303 = 11'h512 == _T_12323 ? mem_1298 : _GEN_1302;
  assign _GEN_1304 = 11'h513 == _T_12323 ? mem_1299 : _GEN_1303;
  assign _GEN_1305 = 11'h514 == _T_12323 ? mem_1300 : _GEN_1304;
  assign _GEN_1306 = 11'h515 == _T_12323 ? mem_1301 : _GEN_1305;
  assign _GEN_1307 = 11'h516 == _T_12323 ? mem_1302 : _GEN_1306;
  assign _GEN_1308 = 11'h517 == _T_12323 ? mem_1303 : _GEN_1307;
  assign _GEN_1309 = 11'h518 == _T_12323 ? mem_1304 : _GEN_1308;
  assign _GEN_1310 = 11'h519 == _T_12323 ? mem_1305 : _GEN_1309;
  assign _GEN_1311 = 11'h51a == _T_12323 ? mem_1306 : _GEN_1310;
  assign _GEN_1312 = 11'h51b == _T_12323 ? mem_1307 : _GEN_1311;
  assign _GEN_1313 = 11'h51c == _T_12323 ? mem_1308 : _GEN_1312;
  assign _GEN_1314 = 11'h51d == _T_12323 ? mem_1309 : _GEN_1313;
  assign _GEN_1315 = 11'h51e == _T_12323 ? mem_1310 : _GEN_1314;
  assign _GEN_1316 = 11'h51f == _T_12323 ? mem_1311 : _GEN_1315;
  assign _GEN_1317 = 11'h520 == _T_12323 ? mem_1312 : _GEN_1316;
  assign _GEN_1318 = 11'h521 == _T_12323 ? mem_1313 : _GEN_1317;
  assign _GEN_1319 = 11'h522 == _T_12323 ? mem_1314 : _GEN_1318;
  assign _GEN_1320 = 11'h523 == _T_12323 ? mem_1315 : _GEN_1319;
  assign _GEN_1321 = 11'h524 == _T_12323 ? mem_1316 : _GEN_1320;
  assign _GEN_1322 = 11'h525 == _T_12323 ? mem_1317 : _GEN_1321;
  assign _GEN_1323 = 11'h526 == _T_12323 ? mem_1318 : _GEN_1322;
  assign _GEN_1324 = 11'h527 == _T_12323 ? mem_1319 : _GEN_1323;
  assign _GEN_1325 = 11'h528 == _T_12323 ? mem_1320 : _GEN_1324;
  assign _GEN_1326 = 11'h529 == _T_12323 ? mem_1321 : _GEN_1325;
  assign _GEN_1327 = 11'h52a == _T_12323 ? mem_1322 : _GEN_1326;
  assign _GEN_1328 = 11'h52b == _T_12323 ? mem_1323 : _GEN_1327;
  assign _GEN_1329 = 11'h52c == _T_12323 ? mem_1324 : _GEN_1328;
  assign _GEN_1330 = 11'h52d == _T_12323 ? mem_1325 : _GEN_1329;
  assign _GEN_1331 = 11'h52e == _T_12323 ? mem_1326 : _GEN_1330;
  assign _GEN_1332 = 11'h52f == _T_12323 ? mem_1327 : _GEN_1331;
  assign _GEN_1333 = 11'h530 == _T_12323 ? mem_1328 : _GEN_1332;
  assign _GEN_1334 = 11'h531 == _T_12323 ? mem_1329 : _GEN_1333;
  assign _GEN_1335 = 11'h532 == _T_12323 ? mem_1330 : _GEN_1334;
  assign _GEN_1336 = 11'h533 == _T_12323 ? mem_1331 : _GEN_1335;
  assign _GEN_1337 = 11'h534 == _T_12323 ? mem_1332 : _GEN_1336;
  assign _GEN_1338 = 11'h535 == _T_12323 ? mem_1333 : _GEN_1337;
  assign _GEN_1339 = 11'h536 == _T_12323 ? mem_1334 : _GEN_1338;
  assign _GEN_1340 = 11'h537 == _T_12323 ? mem_1335 : _GEN_1339;
  assign _GEN_1341 = 11'h538 == _T_12323 ? mem_1336 : _GEN_1340;
  assign _GEN_1342 = 11'h539 == _T_12323 ? mem_1337 : _GEN_1341;
  assign _GEN_1343 = 11'h53a == _T_12323 ? mem_1338 : _GEN_1342;
  assign _GEN_1344 = 11'h53b == _T_12323 ? mem_1339 : _GEN_1343;
  assign _GEN_1345 = 11'h53c == _T_12323 ? mem_1340 : _GEN_1344;
  assign _GEN_1346 = 11'h53d == _T_12323 ? mem_1341 : _GEN_1345;
  assign _GEN_1347 = 11'h53e == _T_12323 ? mem_1342 : _GEN_1346;
  assign _GEN_1348 = 11'h53f == _T_12323 ? mem_1343 : _GEN_1347;
  assign _GEN_1349 = 11'h540 == _T_12323 ? mem_1344 : _GEN_1348;
  assign _GEN_1350 = 11'h541 == _T_12323 ? mem_1345 : _GEN_1349;
  assign _GEN_1351 = 11'h542 == _T_12323 ? mem_1346 : _GEN_1350;
  assign _GEN_1352 = 11'h543 == _T_12323 ? mem_1347 : _GEN_1351;
  assign _GEN_1353 = 11'h544 == _T_12323 ? mem_1348 : _GEN_1352;
  assign _GEN_1354 = 11'h545 == _T_12323 ? mem_1349 : _GEN_1353;
  assign _GEN_1355 = 11'h546 == _T_12323 ? mem_1350 : _GEN_1354;
  assign _GEN_1356 = 11'h547 == _T_12323 ? mem_1351 : _GEN_1355;
  assign _GEN_1357 = 11'h548 == _T_12323 ? mem_1352 : _GEN_1356;
  assign _GEN_1358 = 11'h549 == _T_12323 ? mem_1353 : _GEN_1357;
  assign _GEN_1359 = 11'h54a == _T_12323 ? mem_1354 : _GEN_1358;
  assign _GEN_1360 = 11'h54b == _T_12323 ? mem_1355 : _GEN_1359;
  assign _GEN_1361 = 11'h54c == _T_12323 ? mem_1356 : _GEN_1360;
  assign _GEN_1362 = 11'h54d == _T_12323 ? mem_1357 : _GEN_1361;
  assign _GEN_1363 = 11'h54e == _T_12323 ? mem_1358 : _GEN_1362;
  assign _GEN_1364 = 11'h54f == _T_12323 ? mem_1359 : _GEN_1363;
  assign _GEN_1365 = 11'h550 == _T_12323 ? mem_1360 : _GEN_1364;
  assign _GEN_1366 = 11'h551 == _T_12323 ? mem_1361 : _GEN_1365;
  assign _GEN_1367 = 11'h552 == _T_12323 ? mem_1362 : _GEN_1366;
  assign _GEN_1368 = 11'h553 == _T_12323 ? mem_1363 : _GEN_1367;
  assign _GEN_1369 = 11'h554 == _T_12323 ? mem_1364 : _GEN_1368;
  assign _GEN_1370 = 11'h555 == _T_12323 ? mem_1365 : _GEN_1369;
  assign _GEN_1371 = 11'h556 == _T_12323 ? mem_1366 : _GEN_1370;
  assign _GEN_1372 = 11'h557 == _T_12323 ? mem_1367 : _GEN_1371;
  assign _GEN_1373 = 11'h558 == _T_12323 ? mem_1368 : _GEN_1372;
  assign _GEN_1374 = 11'h559 == _T_12323 ? mem_1369 : _GEN_1373;
  assign _GEN_1375 = 11'h55a == _T_12323 ? mem_1370 : _GEN_1374;
  assign _GEN_1376 = 11'h55b == _T_12323 ? mem_1371 : _GEN_1375;
  assign _GEN_1377 = 11'h55c == _T_12323 ? mem_1372 : _GEN_1376;
  assign _GEN_1378 = 11'h55d == _T_12323 ? mem_1373 : _GEN_1377;
  assign _GEN_1379 = 11'h55e == _T_12323 ? mem_1374 : _GEN_1378;
  assign _GEN_1380 = 11'h55f == _T_12323 ? mem_1375 : _GEN_1379;
  assign _GEN_1381 = 11'h560 == _T_12323 ? mem_1376 : _GEN_1380;
  assign _GEN_1382 = 11'h561 == _T_12323 ? mem_1377 : _GEN_1381;
  assign _GEN_1383 = 11'h562 == _T_12323 ? mem_1378 : _GEN_1382;
  assign _GEN_1384 = 11'h563 == _T_12323 ? mem_1379 : _GEN_1383;
  assign _GEN_1385 = 11'h564 == _T_12323 ? mem_1380 : _GEN_1384;
  assign _GEN_1386 = 11'h565 == _T_12323 ? mem_1381 : _GEN_1385;
  assign _GEN_1387 = 11'h566 == _T_12323 ? mem_1382 : _GEN_1386;
  assign _GEN_1388 = 11'h567 == _T_12323 ? mem_1383 : _GEN_1387;
  assign _GEN_1389 = 11'h568 == _T_12323 ? mem_1384 : _GEN_1388;
  assign _GEN_1390 = 11'h569 == _T_12323 ? mem_1385 : _GEN_1389;
  assign _GEN_1391 = 11'h56a == _T_12323 ? mem_1386 : _GEN_1390;
  assign _GEN_1392 = 11'h56b == _T_12323 ? mem_1387 : _GEN_1391;
  assign _GEN_1393 = 11'h56c == _T_12323 ? mem_1388 : _GEN_1392;
  assign _GEN_1394 = 11'h56d == _T_12323 ? mem_1389 : _GEN_1393;
  assign _GEN_1395 = 11'h56e == _T_12323 ? mem_1390 : _GEN_1394;
  assign _GEN_1396 = 11'h56f == _T_12323 ? mem_1391 : _GEN_1395;
  assign _GEN_1397 = 11'h570 == _T_12323 ? mem_1392 : _GEN_1396;
  assign _GEN_1398 = 11'h571 == _T_12323 ? mem_1393 : _GEN_1397;
  assign _GEN_1399 = 11'h572 == _T_12323 ? mem_1394 : _GEN_1398;
  assign _GEN_1400 = 11'h573 == _T_12323 ? mem_1395 : _GEN_1399;
  assign _GEN_1401 = 11'h574 == _T_12323 ? mem_1396 : _GEN_1400;
  assign _GEN_1402 = 11'h575 == _T_12323 ? mem_1397 : _GEN_1401;
  assign _GEN_1403 = 11'h576 == _T_12323 ? mem_1398 : _GEN_1402;
  assign _GEN_1404 = 11'h577 == _T_12323 ? mem_1399 : _GEN_1403;
  assign _GEN_1405 = 11'h578 == _T_12323 ? mem_1400 : _GEN_1404;
  assign _GEN_1406 = 11'h579 == _T_12323 ? mem_1401 : _GEN_1405;
  assign _GEN_1407 = 11'h57a == _T_12323 ? mem_1402 : _GEN_1406;
  assign _GEN_1408 = 11'h57b == _T_12323 ? mem_1403 : _GEN_1407;
  assign _GEN_1409 = 11'h57c == _T_12323 ? mem_1404 : _GEN_1408;
  assign _GEN_1410 = 11'h57d == _T_12323 ? mem_1405 : _GEN_1409;
  assign _GEN_1411 = 11'h57e == _T_12323 ? mem_1406 : _GEN_1410;
  assign _GEN_1412 = 11'h57f == _T_12323 ? mem_1407 : _GEN_1411;
  assign _GEN_1413 = 11'h580 == _T_12323 ? mem_1408 : _GEN_1412;
  assign _GEN_1414 = 11'h581 == _T_12323 ? mem_1409 : _GEN_1413;
  assign _GEN_1415 = 11'h582 == _T_12323 ? mem_1410 : _GEN_1414;
  assign _GEN_1416 = 11'h583 == _T_12323 ? mem_1411 : _GEN_1415;
  assign _GEN_1417 = 11'h584 == _T_12323 ? mem_1412 : _GEN_1416;
  assign _GEN_1418 = 11'h585 == _T_12323 ? mem_1413 : _GEN_1417;
  assign _GEN_1419 = 11'h586 == _T_12323 ? mem_1414 : _GEN_1418;
  assign _GEN_1420 = 11'h587 == _T_12323 ? mem_1415 : _GEN_1419;
  assign _GEN_1421 = 11'h588 == _T_12323 ? mem_1416 : _GEN_1420;
  assign _GEN_1422 = 11'h589 == _T_12323 ? mem_1417 : _GEN_1421;
  assign _GEN_1423 = 11'h58a == _T_12323 ? mem_1418 : _GEN_1422;
  assign _GEN_1424 = 11'h58b == _T_12323 ? mem_1419 : _GEN_1423;
  assign _GEN_1425 = 11'h58c == _T_12323 ? mem_1420 : _GEN_1424;
  assign _GEN_1426 = 11'h58d == _T_12323 ? mem_1421 : _GEN_1425;
  assign _GEN_1427 = 11'h58e == _T_12323 ? mem_1422 : _GEN_1426;
  assign _GEN_1428 = 11'h58f == _T_12323 ? mem_1423 : _GEN_1427;
  assign _GEN_1429 = 11'h590 == _T_12323 ? mem_1424 : _GEN_1428;
  assign _GEN_1430 = 11'h591 == _T_12323 ? mem_1425 : _GEN_1429;
  assign _GEN_1431 = 11'h592 == _T_12323 ? mem_1426 : _GEN_1430;
  assign _GEN_1432 = 11'h593 == _T_12323 ? mem_1427 : _GEN_1431;
  assign _GEN_1433 = 11'h594 == _T_12323 ? mem_1428 : _GEN_1432;
  assign _GEN_1434 = 11'h595 == _T_12323 ? mem_1429 : _GEN_1433;
  assign _GEN_1435 = 11'h596 == _T_12323 ? mem_1430 : _GEN_1434;
  assign _GEN_1436 = 11'h597 == _T_12323 ? mem_1431 : _GEN_1435;
  assign _GEN_1437 = 11'h598 == _T_12323 ? mem_1432 : _GEN_1436;
  assign _GEN_1438 = 11'h599 == _T_12323 ? mem_1433 : _GEN_1437;
  assign _GEN_1439 = 11'h59a == _T_12323 ? mem_1434 : _GEN_1438;
  assign _GEN_1440 = 11'h59b == _T_12323 ? mem_1435 : _GEN_1439;
  assign _GEN_1441 = 11'h59c == _T_12323 ? mem_1436 : _GEN_1440;
  assign _GEN_1442 = 11'h59d == _T_12323 ? mem_1437 : _GEN_1441;
  assign _GEN_1443 = 11'h59e == _T_12323 ? mem_1438 : _GEN_1442;
  assign _GEN_1444 = 11'h59f == _T_12323 ? mem_1439 : _GEN_1443;
  assign _GEN_1445 = 11'h5a0 == _T_12323 ? mem_1440 : _GEN_1444;
  assign _GEN_1446 = 11'h5a1 == _T_12323 ? mem_1441 : _GEN_1445;
  assign _GEN_1447 = 11'h5a2 == _T_12323 ? mem_1442 : _GEN_1446;
  assign _GEN_1448 = 11'h5a3 == _T_12323 ? mem_1443 : _GEN_1447;
  assign _GEN_1449 = 11'h5a4 == _T_12323 ? mem_1444 : _GEN_1448;
  assign _GEN_1450 = 11'h5a5 == _T_12323 ? mem_1445 : _GEN_1449;
  assign _GEN_1451 = 11'h5a6 == _T_12323 ? mem_1446 : _GEN_1450;
  assign _GEN_1452 = 11'h5a7 == _T_12323 ? mem_1447 : _GEN_1451;
  assign _GEN_1453 = 11'h5a8 == _T_12323 ? mem_1448 : _GEN_1452;
  assign _GEN_1454 = 11'h5a9 == _T_12323 ? mem_1449 : _GEN_1453;
  assign _GEN_1455 = 11'h5aa == _T_12323 ? mem_1450 : _GEN_1454;
  assign _GEN_1456 = 11'h5ab == _T_12323 ? mem_1451 : _GEN_1455;
  assign _GEN_1457 = 11'h5ac == _T_12323 ? mem_1452 : _GEN_1456;
  assign _GEN_1458 = 11'h5ad == _T_12323 ? mem_1453 : _GEN_1457;
  assign _GEN_1459 = 11'h5ae == _T_12323 ? mem_1454 : _GEN_1458;
  assign _GEN_1460 = 11'h5af == _T_12323 ? mem_1455 : _GEN_1459;
  assign _GEN_1461 = 11'h5b0 == _T_12323 ? mem_1456 : _GEN_1460;
  assign _GEN_1462 = 11'h5b1 == _T_12323 ? mem_1457 : _GEN_1461;
  assign _GEN_1463 = 11'h5b2 == _T_12323 ? mem_1458 : _GEN_1462;
  assign _GEN_1464 = 11'h5b3 == _T_12323 ? mem_1459 : _GEN_1463;
  assign _GEN_1465 = 11'h5b4 == _T_12323 ? mem_1460 : _GEN_1464;
  assign _GEN_1466 = 11'h5b5 == _T_12323 ? mem_1461 : _GEN_1465;
  assign _GEN_1467 = 11'h5b6 == _T_12323 ? mem_1462 : _GEN_1466;
  assign _GEN_1468 = 11'h5b7 == _T_12323 ? mem_1463 : _GEN_1467;
  assign _GEN_1469 = 11'h5b8 == _T_12323 ? mem_1464 : _GEN_1468;
  assign _GEN_1470 = 11'h5b9 == _T_12323 ? mem_1465 : _GEN_1469;
  assign _GEN_1471 = 11'h5ba == _T_12323 ? mem_1466 : _GEN_1470;
  assign _GEN_1472 = 11'h5bb == _T_12323 ? mem_1467 : _GEN_1471;
  assign _GEN_1473 = 11'h5bc == _T_12323 ? mem_1468 : _GEN_1472;
  assign _GEN_1474 = 11'h5bd == _T_12323 ? mem_1469 : _GEN_1473;
  assign _GEN_1475 = 11'h5be == _T_12323 ? mem_1470 : _GEN_1474;
  assign _GEN_1476 = 11'h5bf == _T_12323 ? mem_1471 : _GEN_1475;
  assign _GEN_1477 = 11'h5c0 == _T_12323 ? mem_1472 : _GEN_1476;
  assign _GEN_1478 = 11'h5c1 == _T_12323 ? mem_1473 : _GEN_1477;
  assign _GEN_1479 = 11'h5c2 == _T_12323 ? mem_1474 : _GEN_1478;
  assign _GEN_1480 = 11'h5c3 == _T_12323 ? mem_1475 : _GEN_1479;
  assign _GEN_1481 = 11'h5c4 == _T_12323 ? mem_1476 : _GEN_1480;
  assign _GEN_1482 = 11'h5c5 == _T_12323 ? mem_1477 : _GEN_1481;
  assign _GEN_1483 = 11'h5c6 == _T_12323 ? mem_1478 : _GEN_1482;
  assign _GEN_1484 = 11'h5c7 == _T_12323 ? mem_1479 : _GEN_1483;
  assign _GEN_1485 = 11'h5c8 == _T_12323 ? mem_1480 : _GEN_1484;
  assign _GEN_1486 = 11'h5c9 == _T_12323 ? mem_1481 : _GEN_1485;
  assign _GEN_1487 = 11'h5ca == _T_12323 ? mem_1482 : _GEN_1486;
  assign _GEN_1488 = 11'h5cb == _T_12323 ? mem_1483 : _GEN_1487;
  assign _GEN_1489 = 11'h5cc == _T_12323 ? mem_1484 : _GEN_1488;
  assign _GEN_1490 = 11'h5cd == _T_12323 ? mem_1485 : _GEN_1489;
  assign _GEN_1491 = 11'h5ce == _T_12323 ? mem_1486 : _GEN_1490;
  assign _GEN_1492 = 11'h5cf == _T_12323 ? mem_1487 : _GEN_1491;
  assign _GEN_1493 = 11'h5d0 == _T_12323 ? mem_1488 : _GEN_1492;
  assign _GEN_1494 = 11'h5d1 == _T_12323 ? mem_1489 : _GEN_1493;
  assign _GEN_1495 = 11'h5d2 == _T_12323 ? mem_1490 : _GEN_1494;
  assign _GEN_1496 = 11'h5d3 == _T_12323 ? mem_1491 : _GEN_1495;
  assign _GEN_1497 = 11'h5d4 == _T_12323 ? mem_1492 : _GEN_1496;
  assign _GEN_1498 = 11'h5d5 == _T_12323 ? mem_1493 : _GEN_1497;
  assign _GEN_1499 = 11'h5d6 == _T_12323 ? mem_1494 : _GEN_1498;
  assign _GEN_1500 = 11'h5d7 == _T_12323 ? mem_1495 : _GEN_1499;
  assign _GEN_1501 = 11'h5d8 == _T_12323 ? mem_1496 : _GEN_1500;
  assign _GEN_1502 = 11'h5d9 == _T_12323 ? mem_1497 : _GEN_1501;
  assign _GEN_1503 = 11'h5da == _T_12323 ? mem_1498 : _GEN_1502;
  assign _GEN_1504 = 11'h5db == _T_12323 ? mem_1499 : _GEN_1503;
  assign _GEN_1505 = 11'h5dc == _T_12323 ? mem_1500 : _GEN_1504;
  assign _GEN_1506 = 11'h5dd == _T_12323 ? mem_1501 : _GEN_1505;
  assign _GEN_1507 = 11'h5de == _T_12323 ? mem_1502 : _GEN_1506;
  assign _GEN_1508 = 11'h5df == _T_12323 ? mem_1503 : _GEN_1507;
  assign _GEN_1509 = 11'h5e0 == _T_12323 ? mem_1504 : _GEN_1508;
  assign _GEN_1510 = 11'h5e1 == _T_12323 ? mem_1505 : _GEN_1509;
  assign _GEN_1511 = 11'h5e2 == _T_12323 ? mem_1506 : _GEN_1510;
  assign _GEN_1512 = 11'h5e3 == _T_12323 ? mem_1507 : _GEN_1511;
  assign _GEN_1513 = 11'h5e4 == _T_12323 ? mem_1508 : _GEN_1512;
  assign _GEN_1514 = 11'h5e5 == _T_12323 ? mem_1509 : _GEN_1513;
  assign _GEN_1515 = 11'h5e6 == _T_12323 ? mem_1510 : _GEN_1514;
  assign _GEN_1516 = 11'h5e7 == _T_12323 ? mem_1511 : _GEN_1515;
  assign _GEN_1517 = 11'h5e8 == _T_12323 ? mem_1512 : _GEN_1516;
  assign _GEN_1518 = 11'h5e9 == _T_12323 ? mem_1513 : _GEN_1517;
  assign _GEN_1519 = 11'h5ea == _T_12323 ? mem_1514 : _GEN_1518;
  assign _GEN_1520 = 11'h5eb == _T_12323 ? mem_1515 : _GEN_1519;
  assign _GEN_1521 = 11'h5ec == _T_12323 ? mem_1516 : _GEN_1520;
  assign _GEN_1522 = 11'h5ed == _T_12323 ? mem_1517 : _GEN_1521;
  assign _GEN_1523 = 11'h5ee == _T_12323 ? mem_1518 : _GEN_1522;
  assign _GEN_1524 = 11'h5ef == _T_12323 ? mem_1519 : _GEN_1523;
  assign _GEN_1525 = 11'h5f0 == _T_12323 ? mem_1520 : _GEN_1524;
  assign _GEN_1526 = 11'h5f1 == _T_12323 ? mem_1521 : _GEN_1525;
  assign _GEN_1527 = 11'h5f2 == _T_12323 ? mem_1522 : _GEN_1526;
  assign _GEN_1528 = 11'h5f3 == _T_12323 ? mem_1523 : _GEN_1527;
  assign _GEN_1529 = 11'h5f4 == _T_12323 ? mem_1524 : _GEN_1528;
  assign _GEN_1530 = 11'h5f5 == _T_12323 ? mem_1525 : _GEN_1529;
  assign _GEN_1531 = 11'h5f6 == _T_12323 ? mem_1526 : _GEN_1530;
  assign _GEN_1532 = 11'h5f7 == _T_12323 ? mem_1527 : _GEN_1531;
  assign _GEN_1533 = 11'h5f8 == _T_12323 ? mem_1528 : _GEN_1532;
  assign _GEN_1534 = 11'h5f9 == _T_12323 ? mem_1529 : _GEN_1533;
  assign _GEN_1535 = 11'h5fa == _T_12323 ? mem_1530 : _GEN_1534;
  assign _GEN_1536 = 11'h5fb == _T_12323 ? mem_1531 : _GEN_1535;
  assign _GEN_1537 = 11'h5fc == _T_12323 ? mem_1532 : _GEN_1536;
  assign _GEN_1538 = 11'h5fd == _T_12323 ? mem_1533 : _GEN_1537;
  assign _GEN_1539 = 11'h5fe == _T_12323 ? mem_1534 : _GEN_1538;
  assign _GEN_1540 = 11'h5ff == _T_12323 ? mem_1535 : _GEN_1539;
  assign _GEN_1541 = 11'h600 == _T_12323 ? mem_1536 : _GEN_1540;
  assign _GEN_1542 = 11'h601 == _T_12323 ? mem_1537 : _GEN_1541;
  assign _GEN_1543 = 11'h602 == _T_12323 ? mem_1538 : _GEN_1542;
  assign _GEN_1544 = 11'h603 == _T_12323 ? mem_1539 : _GEN_1543;
  assign _GEN_1545 = 11'h604 == _T_12323 ? mem_1540 : _GEN_1544;
  assign _GEN_1546 = 11'h605 == _T_12323 ? mem_1541 : _GEN_1545;
  assign _GEN_1547 = 11'h606 == _T_12323 ? mem_1542 : _GEN_1546;
  assign _GEN_1548 = 11'h607 == _T_12323 ? mem_1543 : _GEN_1547;
  assign _GEN_1549 = 11'h608 == _T_12323 ? mem_1544 : _GEN_1548;
  assign _GEN_1550 = 11'h609 == _T_12323 ? mem_1545 : _GEN_1549;
  assign _GEN_1551 = 11'h60a == _T_12323 ? mem_1546 : _GEN_1550;
  assign _GEN_1552 = 11'h60b == _T_12323 ? mem_1547 : _GEN_1551;
  assign _GEN_1553 = 11'h60c == _T_12323 ? mem_1548 : _GEN_1552;
  assign _GEN_1554 = 11'h60d == _T_12323 ? mem_1549 : _GEN_1553;
  assign _GEN_1555 = 11'h60e == _T_12323 ? mem_1550 : _GEN_1554;
  assign _GEN_1556 = 11'h60f == _T_12323 ? mem_1551 : _GEN_1555;
  assign _GEN_1557 = 11'h610 == _T_12323 ? mem_1552 : _GEN_1556;
  assign _GEN_1558 = 11'h611 == _T_12323 ? mem_1553 : _GEN_1557;
  assign _GEN_1559 = 11'h612 == _T_12323 ? mem_1554 : _GEN_1558;
  assign _GEN_1560 = 11'h613 == _T_12323 ? mem_1555 : _GEN_1559;
  assign _GEN_1561 = 11'h614 == _T_12323 ? mem_1556 : _GEN_1560;
  assign _GEN_1562 = 11'h615 == _T_12323 ? mem_1557 : _GEN_1561;
  assign _GEN_1563 = 11'h616 == _T_12323 ? mem_1558 : _GEN_1562;
  assign _GEN_1564 = 11'h617 == _T_12323 ? mem_1559 : _GEN_1563;
  assign _GEN_1565 = 11'h618 == _T_12323 ? mem_1560 : _GEN_1564;
  assign _GEN_1566 = 11'h619 == _T_12323 ? mem_1561 : _GEN_1565;
  assign _GEN_1567 = 11'h61a == _T_12323 ? mem_1562 : _GEN_1566;
  assign _GEN_1568 = 11'h61b == _T_12323 ? mem_1563 : _GEN_1567;
  assign _GEN_1569 = 11'h61c == _T_12323 ? mem_1564 : _GEN_1568;
  assign _GEN_1570 = 11'h61d == _T_12323 ? mem_1565 : _GEN_1569;
  assign _GEN_1571 = 11'h61e == _T_12323 ? mem_1566 : _GEN_1570;
  assign _GEN_1572 = 11'h61f == _T_12323 ? mem_1567 : _GEN_1571;
  assign _GEN_1573 = 11'h620 == _T_12323 ? mem_1568 : _GEN_1572;
  assign _GEN_1574 = 11'h621 == _T_12323 ? mem_1569 : _GEN_1573;
  assign _GEN_1575 = 11'h622 == _T_12323 ? mem_1570 : _GEN_1574;
  assign _GEN_1576 = 11'h623 == _T_12323 ? mem_1571 : _GEN_1575;
  assign _GEN_1577 = 11'h624 == _T_12323 ? mem_1572 : _GEN_1576;
  assign _GEN_1578 = 11'h625 == _T_12323 ? mem_1573 : _GEN_1577;
  assign _GEN_1579 = 11'h626 == _T_12323 ? mem_1574 : _GEN_1578;
  assign _GEN_1580 = 11'h627 == _T_12323 ? mem_1575 : _GEN_1579;
  assign _GEN_1581 = 11'h628 == _T_12323 ? mem_1576 : _GEN_1580;
  assign _GEN_1582 = 11'h629 == _T_12323 ? mem_1577 : _GEN_1581;
  assign _GEN_1583 = 11'h62a == _T_12323 ? mem_1578 : _GEN_1582;
  assign _GEN_1584 = 11'h62b == _T_12323 ? mem_1579 : _GEN_1583;
  assign _GEN_1585 = 11'h62c == _T_12323 ? mem_1580 : _GEN_1584;
  assign _GEN_1586 = 11'h62d == _T_12323 ? mem_1581 : _GEN_1585;
  assign _GEN_1587 = 11'h62e == _T_12323 ? mem_1582 : _GEN_1586;
  assign _GEN_1588 = 11'h62f == _T_12323 ? mem_1583 : _GEN_1587;
  assign _GEN_1589 = 11'h630 == _T_12323 ? mem_1584 : _GEN_1588;
  assign _GEN_1590 = 11'h631 == _T_12323 ? mem_1585 : _GEN_1589;
  assign _GEN_1591 = 11'h632 == _T_12323 ? mem_1586 : _GEN_1590;
  assign _GEN_1592 = 11'h633 == _T_12323 ? mem_1587 : _GEN_1591;
  assign _GEN_1593 = 11'h634 == _T_12323 ? mem_1588 : _GEN_1592;
  assign _GEN_1594 = 11'h635 == _T_12323 ? mem_1589 : _GEN_1593;
  assign _GEN_1595 = 11'h636 == _T_12323 ? mem_1590 : _GEN_1594;
  assign _GEN_1596 = 11'h637 == _T_12323 ? mem_1591 : _GEN_1595;
  assign _GEN_1597 = 11'h638 == _T_12323 ? mem_1592 : _GEN_1596;
  assign _GEN_1598 = 11'h639 == _T_12323 ? mem_1593 : _GEN_1597;
  assign _GEN_1599 = 11'h63a == _T_12323 ? mem_1594 : _GEN_1598;
  assign _GEN_1600 = 11'h63b == _T_12323 ? mem_1595 : _GEN_1599;
  assign _GEN_1601 = 11'h63c == _T_12323 ? mem_1596 : _GEN_1600;
  assign _GEN_1602 = 11'h63d == _T_12323 ? mem_1597 : _GEN_1601;
  assign _GEN_1603 = 11'h63e == _T_12323 ? mem_1598 : _GEN_1602;
  assign _GEN_1604 = 11'h63f == _T_12323 ? mem_1599 : _GEN_1603;
  assign _GEN_1605 = 11'h640 == _T_12323 ? mem_1600 : _GEN_1604;
  assign _GEN_1606 = 11'h641 == _T_12323 ? mem_1601 : _GEN_1605;
  assign _GEN_1607 = 11'h642 == _T_12323 ? mem_1602 : _GEN_1606;
  assign _GEN_1608 = 11'h643 == _T_12323 ? mem_1603 : _GEN_1607;
  assign _GEN_1609 = 11'h644 == _T_12323 ? mem_1604 : _GEN_1608;
  assign _GEN_1610 = 11'h645 == _T_12323 ? mem_1605 : _GEN_1609;
  assign _GEN_1611 = 11'h646 == _T_12323 ? mem_1606 : _GEN_1610;
  assign _GEN_1612 = 11'h647 == _T_12323 ? mem_1607 : _GEN_1611;
  assign _GEN_1613 = 11'h648 == _T_12323 ? mem_1608 : _GEN_1612;
  assign _GEN_1614 = 11'h649 == _T_12323 ? mem_1609 : _GEN_1613;
  assign _GEN_1615 = 11'h64a == _T_12323 ? mem_1610 : _GEN_1614;
  assign _GEN_1616 = 11'h64b == _T_12323 ? mem_1611 : _GEN_1615;
  assign _GEN_1617 = 11'h64c == _T_12323 ? mem_1612 : _GEN_1616;
  assign _GEN_1618 = 11'h64d == _T_12323 ? mem_1613 : _GEN_1617;
  assign _GEN_1619 = 11'h64e == _T_12323 ? mem_1614 : _GEN_1618;
  assign _GEN_1620 = 11'h64f == _T_12323 ? mem_1615 : _GEN_1619;
  assign _GEN_1621 = 11'h650 == _T_12323 ? mem_1616 : _GEN_1620;
  assign _GEN_1622 = 11'h651 == _T_12323 ? mem_1617 : _GEN_1621;
  assign _GEN_1623 = 11'h652 == _T_12323 ? mem_1618 : _GEN_1622;
  assign _GEN_1624 = 11'h653 == _T_12323 ? mem_1619 : _GEN_1623;
  assign _GEN_1625 = 11'h654 == _T_12323 ? mem_1620 : _GEN_1624;
  assign _GEN_1626 = 11'h655 == _T_12323 ? mem_1621 : _GEN_1625;
  assign _GEN_1627 = 11'h656 == _T_12323 ? mem_1622 : _GEN_1626;
  assign _GEN_1628 = 11'h657 == _T_12323 ? mem_1623 : _GEN_1627;
  assign _GEN_1629 = 11'h658 == _T_12323 ? mem_1624 : _GEN_1628;
  assign _GEN_1630 = 11'h659 == _T_12323 ? mem_1625 : _GEN_1629;
  assign _GEN_1631 = 11'h65a == _T_12323 ? mem_1626 : _GEN_1630;
  assign _GEN_1632 = 11'h65b == _T_12323 ? mem_1627 : _GEN_1631;
  assign _GEN_1633 = 11'h65c == _T_12323 ? mem_1628 : _GEN_1632;
  assign _GEN_1634 = 11'h65d == _T_12323 ? mem_1629 : _GEN_1633;
  assign _GEN_1635 = 11'h65e == _T_12323 ? mem_1630 : _GEN_1634;
  assign _GEN_1636 = 11'h65f == _T_12323 ? mem_1631 : _GEN_1635;
  assign _GEN_1637 = 11'h660 == _T_12323 ? mem_1632 : _GEN_1636;
  assign _GEN_1638 = 11'h661 == _T_12323 ? mem_1633 : _GEN_1637;
  assign _GEN_1639 = 11'h662 == _T_12323 ? mem_1634 : _GEN_1638;
  assign _GEN_1640 = 11'h663 == _T_12323 ? mem_1635 : _GEN_1639;
  assign _GEN_1641 = 11'h664 == _T_12323 ? mem_1636 : _GEN_1640;
  assign _GEN_1642 = 11'h665 == _T_12323 ? mem_1637 : _GEN_1641;
  assign _GEN_1643 = 11'h666 == _T_12323 ? mem_1638 : _GEN_1642;
  assign _GEN_1644 = 11'h667 == _T_12323 ? mem_1639 : _GEN_1643;
  assign _GEN_1645 = 11'h668 == _T_12323 ? mem_1640 : _GEN_1644;
  assign _GEN_1646 = 11'h669 == _T_12323 ? mem_1641 : _GEN_1645;
  assign _GEN_1647 = 11'h66a == _T_12323 ? mem_1642 : _GEN_1646;
  assign _GEN_1648 = 11'h66b == _T_12323 ? mem_1643 : _GEN_1647;
  assign _GEN_1649 = 11'h66c == _T_12323 ? mem_1644 : _GEN_1648;
  assign _GEN_1650 = 11'h66d == _T_12323 ? mem_1645 : _GEN_1649;
  assign _GEN_1651 = 11'h66e == _T_12323 ? mem_1646 : _GEN_1650;
  assign _GEN_1652 = 11'h66f == _T_12323 ? mem_1647 : _GEN_1651;
  assign _GEN_1653 = 11'h670 == _T_12323 ? mem_1648 : _GEN_1652;
  assign _GEN_1654 = 11'h671 == _T_12323 ? mem_1649 : _GEN_1653;
  assign _GEN_1655 = 11'h672 == _T_12323 ? mem_1650 : _GEN_1654;
  assign _GEN_1656 = 11'h673 == _T_12323 ? mem_1651 : _GEN_1655;
  assign _GEN_1657 = 11'h674 == _T_12323 ? mem_1652 : _GEN_1656;
  assign _GEN_1658 = 11'h675 == _T_12323 ? mem_1653 : _GEN_1657;
  assign _GEN_1659 = 11'h676 == _T_12323 ? mem_1654 : _GEN_1658;
  assign _GEN_1660 = 11'h677 == _T_12323 ? mem_1655 : _GEN_1659;
  assign _GEN_1661 = 11'h678 == _T_12323 ? mem_1656 : _GEN_1660;
  assign _GEN_1662 = 11'h679 == _T_12323 ? mem_1657 : _GEN_1661;
  assign _GEN_1663 = 11'h67a == _T_12323 ? mem_1658 : _GEN_1662;
  assign _GEN_1664 = 11'h67b == _T_12323 ? mem_1659 : _GEN_1663;
  assign _GEN_1665 = 11'h67c == _T_12323 ? mem_1660 : _GEN_1664;
  assign _GEN_1666 = 11'h67d == _T_12323 ? mem_1661 : _GEN_1665;
  assign _GEN_1667 = 11'h67e == _T_12323 ? mem_1662 : _GEN_1666;
  assign _GEN_1668 = 11'h67f == _T_12323 ? mem_1663 : _GEN_1667;
  assign _GEN_1669 = 11'h680 == _T_12323 ? mem_1664 : _GEN_1668;
  assign _GEN_1670 = 11'h681 == _T_12323 ? mem_1665 : _GEN_1669;
  assign _GEN_1671 = 11'h682 == _T_12323 ? mem_1666 : _GEN_1670;
  assign _GEN_1672 = 11'h683 == _T_12323 ? mem_1667 : _GEN_1671;
  assign _GEN_1673 = 11'h684 == _T_12323 ? mem_1668 : _GEN_1672;
  assign _GEN_1674 = 11'h685 == _T_12323 ? mem_1669 : _GEN_1673;
  assign _GEN_1675 = 11'h686 == _T_12323 ? mem_1670 : _GEN_1674;
  assign _GEN_1676 = 11'h687 == _T_12323 ? mem_1671 : _GEN_1675;
  assign _GEN_1677 = 11'h688 == _T_12323 ? mem_1672 : _GEN_1676;
  assign _GEN_1678 = 11'h689 == _T_12323 ? mem_1673 : _GEN_1677;
  assign _GEN_1679 = 11'h68a == _T_12323 ? mem_1674 : _GEN_1678;
  assign _GEN_1680 = 11'h68b == _T_12323 ? mem_1675 : _GEN_1679;
  assign _GEN_1681 = 11'h68c == _T_12323 ? mem_1676 : _GEN_1680;
  assign _GEN_1682 = 11'h68d == _T_12323 ? mem_1677 : _GEN_1681;
  assign _GEN_1683 = 11'h68e == _T_12323 ? mem_1678 : _GEN_1682;
  assign _GEN_1684 = 11'h68f == _T_12323 ? mem_1679 : _GEN_1683;
  assign _GEN_1685 = 11'h690 == _T_12323 ? mem_1680 : _GEN_1684;
  assign _GEN_1686 = 11'h691 == _T_12323 ? mem_1681 : _GEN_1685;
  assign _GEN_1687 = 11'h692 == _T_12323 ? mem_1682 : _GEN_1686;
  assign _GEN_1688 = 11'h693 == _T_12323 ? mem_1683 : _GEN_1687;
  assign _GEN_1689 = 11'h694 == _T_12323 ? mem_1684 : _GEN_1688;
  assign _GEN_1690 = 11'h695 == _T_12323 ? mem_1685 : _GEN_1689;
  assign _GEN_1691 = 11'h696 == _T_12323 ? mem_1686 : _GEN_1690;
  assign _GEN_1692 = 11'h697 == _T_12323 ? mem_1687 : _GEN_1691;
  assign _GEN_1693 = 11'h698 == _T_12323 ? mem_1688 : _GEN_1692;
  assign _GEN_1694 = 11'h699 == _T_12323 ? mem_1689 : _GEN_1693;
  assign _GEN_1695 = 11'h69a == _T_12323 ? mem_1690 : _GEN_1694;
  assign _GEN_1696 = 11'h69b == _T_12323 ? mem_1691 : _GEN_1695;
  assign _GEN_1697 = 11'h69c == _T_12323 ? mem_1692 : _GEN_1696;
  assign _GEN_1698 = 11'h69d == _T_12323 ? mem_1693 : _GEN_1697;
  assign _GEN_1699 = 11'h69e == _T_12323 ? mem_1694 : _GEN_1698;
  assign _GEN_1700 = 11'h69f == _T_12323 ? mem_1695 : _GEN_1699;
  assign _GEN_1701 = 11'h6a0 == _T_12323 ? mem_1696 : _GEN_1700;
  assign _GEN_1702 = 11'h6a1 == _T_12323 ? mem_1697 : _GEN_1701;
  assign _GEN_1703 = 11'h6a2 == _T_12323 ? mem_1698 : _GEN_1702;
  assign _GEN_1704 = 11'h6a3 == _T_12323 ? mem_1699 : _GEN_1703;
  assign _GEN_1705 = 11'h6a4 == _T_12323 ? mem_1700 : _GEN_1704;
  assign _GEN_1706 = 11'h6a5 == _T_12323 ? mem_1701 : _GEN_1705;
  assign _GEN_1707 = 11'h6a6 == _T_12323 ? mem_1702 : _GEN_1706;
  assign _GEN_1708 = 11'h6a7 == _T_12323 ? mem_1703 : _GEN_1707;
  assign _GEN_1709 = 11'h6a8 == _T_12323 ? mem_1704 : _GEN_1708;
  assign _GEN_1710 = 11'h6a9 == _T_12323 ? mem_1705 : _GEN_1709;
  assign _GEN_1711 = 11'h6aa == _T_12323 ? mem_1706 : _GEN_1710;
  assign _GEN_1712 = 11'h6ab == _T_12323 ? mem_1707 : _GEN_1711;
  assign _GEN_1713 = 11'h6ac == _T_12323 ? mem_1708 : _GEN_1712;
  assign _GEN_1714 = 11'h6ad == _T_12323 ? mem_1709 : _GEN_1713;
  assign _GEN_1715 = 11'h6ae == _T_12323 ? mem_1710 : _GEN_1714;
  assign _GEN_1716 = 11'h6af == _T_12323 ? mem_1711 : _GEN_1715;
  assign _GEN_1717 = 11'h6b0 == _T_12323 ? mem_1712 : _GEN_1716;
  assign _GEN_1718 = 11'h6b1 == _T_12323 ? mem_1713 : _GEN_1717;
  assign _GEN_1719 = 11'h6b2 == _T_12323 ? mem_1714 : _GEN_1718;
  assign _GEN_1720 = 11'h6b3 == _T_12323 ? mem_1715 : _GEN_1719;
  assign _GEN_1721 = 11'h6b4 == _T_12323 ? mem_1716 : _GEN_1720;
  assign _GEN_1722 = 11'h6b5 == _T_12323 ? mem_1717 : _GEN_1721;
  assign _GEN_1723 = 11'h6b6 == _T_12323 ? mem_1718 : _GEN_1722;
  assign _GEN_1724 = 11'h6b7 == _T_12323 ? mem_1719 : _GEN_1723;
  assign _GEN_1725 = 11'h6b8 == _T_12323 ? mem_1720 : _GEN_1724;
  assign _GEN_1726 = 11'h6b9 == _T_12323 ? mem_1721 : _GEN_1725;
  assign _GEN_1727 = 11'h6ba == _T_12323 ? mem_1722 : _GEN_1726;
  assign _GEN_1728 = 11'h6bb == _T_12323 ? mem_1723 : _GEN_1727;
  assign _GEN_1729 = 11'h6bc == _T_12323 ? mem_1724 : _GEN_1728;
  assign _GEN_1730 = 11'h6bd == _T_12323 ? mem_1725 : _GEN_1729;
  assign _GEN_1731 = 11'h6be == _T_12323 ? mem_1726 : _GEN_1730;
  assign _GEN_1732 = 11'h6bf == _T_12323 ? mem_1727 : _GEN_1731;
  assign _GEN_1733 = 11'h6c0 == _T_12323 ? mem_1728 : _GEN_1732;
  assign _GEN_1734 = 11'h6c1 == _T_12323 ? mem_1729 : _GEN_1733;
  assign _GEN_1735 = 11'h6c2 == _T_12323 ? mem_1730 : _GEN_1734;
  assign _GEN_1736 = 11'h6c3 == _T_12323 ? mem_1731 : _GEN_1735;
  assign _GEN_1737 = 11'h6c4 == _T_12323 ? mem_1732 : _GEN_1736;
  assign _GEN_1738 = 11'h6c5 == _T_12323 ? mem_1733 : _GEN_1737;
  assign _GEN_1739 = 11'h6c6 == _T_12323 ? mem_1734 : _GEN_1738;
  assign _GEN_1740 = 11'h6c7 == _T_12323 ? mem_1735 : _GEN_1739;
  assign _GEN_1741 = 11'h6c8 == _T_12323 ? mem_1736 : _GEN_1740;
  assign _GEN_1742 = 11'h6c9 == _T_12323 ? mem_1737 : _GEN_1741;
  assign _GEN_1743 = 11'h6ca == _T_12323 ? mem_1738 : _GEN_1742;
  assign _GEN_1744 = 11'h6cb == _T_12323 ? mem_1739 : _GEN_1743;
  assign _GEN_1745 = 11'h6cc == _T_12323 ? mem_1740 : _GEN_1744;
  assign _GEN_1746 = 11'h6cd == _T_12323 ? mem_1741 : _GEN_1745;
  assign _GEN_1747 = 11'h6ce == _T_12323 ? mem_1742 : _GEN_1746;
  assign _GEN_1748 = 11'h6cf == _T_12323 ? mem_1743 : _GEN_1747;
  assign _GEN_1749 = 11'h6d0 == _T_12323 ? mem_1744 : _GEN_1748;
  assign _GEN_1750 = 11'h6d1 == _T_12323 ? mem_1745 : _GEN_1749;
  assign _GEN_1751 = 11'h6d2 == _T_12323 ? mem_1746 : _GEN_1750;
  assign _GEN_1752 = 11'h6d3 == _T_12323 ? mem_1747 : _GEN_1751;
  assign _GEN_1753 = 11'h6d4 == _T_12323 ? mem_1748 : _GEN_1752;
  assign _GEN_1754 = 11'h6d5 == _T_12323 ? mem_1749 : _GEN_1753;
  assign _GEN_1755 = 11'h6d6 == _T_12323 ? mem_1750 : _GEN_1754;
  assign _GEN_1756 = 11'h6d7 == _T_12323 ? mem_1751 : _GEN_1755;
  assign _GEN_1757 = 11'h6d8 == _T_12323 ? mem_1752 : _GEN_1756;
  assign _GEN_1758 = 11'h6d9 == _T_12323 ? mem_1753 : _GEN_1757;
  assign _GEN_1759 = 11'h6da == _T_12323 ? mem_1754 : _GEN_1758;
  assign _GEN_1760 = 11'h6db == _T_12323 ? mem_1755 : _GEN_1759;
  assign _GEN_1761 = 11'h6dc == _T_12323 ? mem_1756 : _GEN_1760;
  assign _GEN_1762 = 11'h6dd == _T_12323 ? mem_1757 : _GEN_1761;
  assign _GEN_1763 = 11'h6de == _T_12323 ? mem_1758 : _GEN_1762;
  assign _GEN_1764 = 11'h6df == _T_12323 ? mem_1759 : _GEN_1763;
  assign _GEN_1765 = 11'h6e0 == _T_12323 ? mem_1760 : _GEN_1764;
  assign _GEN_1766 = 11'h6e1 == _T_12323 ? mem_1761 : _GEN_1765;
  assign _GEN_1767 = 11'h6e2 == _T_12323 ? mem_1762 : _GEN_1766;
  assign _GEN_1768 = 11'h6e3 == _T_12323 ? mem_1763 : _GEN_1767;
  assign _GEN_1769 = 11'h6e4 == _T_12323 ? mem_1764 : _GEN_1768;
  assign _GEN_1770 = 11'h6e5 == _T_12323 ? mem_1765 : _GEN_1769;
  assign _GEN_1771 = 11'h6e6 == _T_12323 ? mem_1766 : _GEN_1770;
  assign _GEN_1772 = 11'h6e7 == _T_12323 ? mem_1767 : _GEN_1771;
  assign _GEN_1773 = 11'h6e8 == _T_12323 ? mem_1768 : _GEN_1772;
  assign _GEN_1774 = 11'h6e9 == _T_12323 ? mem_1769 : _GEN_1773;
  assign _GEN_1775 = 11'h6ea == _T_12323 ? mem_1770 : _GEN_1774;
  assign _GEN_1776 = 11'h6eb == _T_12323 ? mem_1771 : _GEN_1775;
  assign _GEN_1777 = 11'h6ec == _T_12323 ? mem_1772 : _GEN_1776;
  assign _GEN_1778 = 11'h6ed == _T_12323 ? mem_1773 : _GEN_1777;
  assign _GEN_1779 = 11'h6ee == _T_12323 ? mem_1774 : _GEN_1778;
  assign _GEN_1780 = 11'h6ef == _T_12323 ? mem_1775 : _GEN_1779;
  assign _GEN_1781 = 11'h6f0 == _T_12323 ? mem_1776 : _GEN_1780;
  assign _GEN_1782 = 11'h6f1 == _T_12323 ? mem_1777 : _GEN_1781;
  assign _GEN_1783 = 11'h6f2 == _T_12323 ? mem_1778 : _GEN_1782;
  assign _GEN_1784 = 11'h6f3 == _T_12323 ? mem_1779 : _GEN_1783;
  assign _GEN_1785 = 11'h6f4 == _T_12323 ? mem_1780 : _GEN_1784;
  assign _GEN_1786 = 11'h6f5 == _T_12323 ? mem_1781 : _GEN_1785;
  assign _GEN_1787 = 11'h6f6 == _T_12323 ? mem_1782 : _GEN_1786;
  assign _GEN_1788 = 11'h6f7 == _T_12323 ? mem_1783 : _GEN_1787;
  assign _GEN_1789 = 11'h6f8 == _T_12323 ? mem_1784 : _GEN_1788;
  assign _GEN_1790 = 11'h6f9 == _T_12323 ? mem_1785 : _GEN_1789;
  assign _GEN_1791 = 11'h6fa == _T_12323 ? mem_1786 : _GEN_1790;
  assign _GEN_1792 = 11'h6fb == _T_12323 ? mem_1787 : _GEN_1791;
  assign _GEN_1793 = 11'h6fc == _T_12323 ? mem_1788 : _GEN_1792;
  assign _GEN_1794 = 11'h6fd == _T_12323 ? mem_1789 : _GEN_1793;
  assign _GEN_1795 = 11'h6fe == _T_12323 ? mem_1790 : _GEN_1794;
  assign _GEN_1796 = 11'h6ff == _T_12323 ? mem_1791 : _GEN_1795;
  assign _GEN_1797 = 11'h700 == _T_12323 ? mem_1792 : _GEN_1796;
  assign _GEN_1798 = 11'h701 == _T_12323 ? mem_1793 : _GEN_1797;
  assign _GEN_1799 = 11'h702 == _T_12323 ? mem_1794 : _GEN_1798;
  assign _GEN_1800 = 11'h703 == _T_12323 ? mem_1795 : _GEN_1799;
  assign _GEN_1801 = 11'h704 == _T_12323 ? mem_1796 : _GEN_1800;
  assign _GEN_1802 = 11'h705 == _T_12323 ? mem_1797 : _GEN_1801;
  assign _GEN_1803 = 11'h706 == _T_12323 ? mem_1798 : _GEN_1802;
  assign _GEN_1804 = 11'h707 == _T_12323 ? mem_1799 : _GEN_1803;
  assign _GEN_1805 = 11'h708 == _T_12323 ? mem_1800 : _GEN_1804;
  assign _GEN_1806 = 11'h709 == _T_12323 ? mem_1801 : _GEN_1805;
  assign _GEN_1807 = 11'h70a == _T_12323 ? mem_1802 : _GEN_1806;
  assign _GEN_1808 = 11'h70b == _T_12323 ? mem_1803 : _GEN_1807;
  assign _GEN_1809 = 11'h70c == _T_12323 ? mem_1804 : _GEN_1808;
  assign _GEN_1810 = 11'h70d == _T_12323 ? mem_1805 : _GEN_1809;
  assign _GEN_1811 = 11'h70e == _T_12323 ? mem_1806 : _GEN_1810;
  assign _GEN_1812 = 11'h70f == _T_12323 ? mem_1807 : _GEN_1811;
  assign _GEN_1813 = 11'h710 == _T_12323 ? mem_1808 : _GEN_1812;
  assign _GEN_1814 = 11'h711 == _T_12323 ? mem_1809 : _GEN_1813;
  assign _GEN_1815 = 11'h712 == _T_12323 ? mem_1810 : _GEN_1814;
  assign _GEN_1816 = 11'h713 == _T_12323 ? mem_1811 : _GEN_1815;
  assign _GEN_1817 = 11'h714 == _T_12323 ? mem_1812 : _GEN_1816;
  assign _GEN_1818 = 11'h715 == _T_12323 ? mem_1813 : _GEN_1817;
  assign _GEN_1819 = 11'h716 == _T_12323 ? mem_1814 : _GEN_1818;
  assign _GEN_1820 = 11'h717 == _T_12323 ? mem_1815 : _GEN_1819;
  assign _GEN_1821 = 11'h718 == _T_12323 ? mem_1816 : _GEN_1820;
  assign _GEN_1822 = 11'h719 == _T_12323 ? mem_1817 : _GEN_1821;
  assign _GEN_1823 = 11'h71a == _T_12323 ? mem_1818 : _GEN_1822;
  assign _GEN_1824 = 11'h71b == _T_12323 ? mem_1819 : _GEN_1823;
  assign _GEN_1825 = 11'h71c == _T_12323 ? mem_1820 : _GEN_1824;
  assign _GEN_1826 = 11'h71d == _T_12323 ? mem_1821 : _GEN_1825;
  assign _GEN_1827 = 11'h71e == _T_12323 ? mem_1822 : _GEN_1826;
  assign _GEN_1828 = 11'h71f == _T_12323 ? mem_1823 : _GEN_1827;
  assign _GEN_1829 = 11'h720 == _T_12323 ? mem_1824 : _GEN_1828;
  assign _GEN_1830 = 11'h721 == _T_12323 ? mem_1825 : _GEN_1829;
  assign _GEN_1831 = 11'h722 == _T_12323 ? mem_1826 : _GEN_1830;
  assign _GEN_1832 = 11'h723 == _T_12323 ? mem_1827 : _GEN_1831;
  assign _GEN_1833 = 11'h724 == _T_12323 ? mem_1828 : _GEN_1832;
  assign _GEN_1834 = 11'h725 == _T_12323 ? mem_1829 : _GEN_1833;
  assign _GEN_1835 = 11'h726 == _T_12323 ? mem_1830 : _GEN_1834;
  assign _GEN_1836 = 11'h727 == _T_12323 ? mem_1831 : _GEN_1835;
  assign _GEN_1837 = 11'h728 == _T_12323 ? mem_1832 : _GEN_1836;
  assign _GEN_1838 = 11'h729 == _T_12323 ? mem_1833 : _GEN_1837;
  assign _GEN_1839 = 11'h72a == _T_12323 ? mem_1834 : _GEN_1838;
  assign _GEN_1840 = 11'h72b == _T_12323 ? mem_1835 : _GEN_1839;
  assign _GEN_1841 = 11'h72c == _T_12323 ? mem_1836 : _GEN_1840;
  assign _GEN_1842 = 11'h72d == _T_12323 ? mem_1837 : _GEN_1841;
  assign _GEN_1843 = 11'h72e == _T_12323 ? mem_1838 : _GEN_1842;
  assign _GEN_1844 = 11'h72f == _T_12323 ? mem_1839 : _GEN_1843;
  assign _GEN_1845 = 11'h730 == _T_12323 ? mem_1840 : _GEN_1844;
  assign _GEN_1846 = 11'h731 == _T_12323 ? mem_1841 : _GEN_1845;
  assign _GEN_1847 = 11'h732 == _T_12323 ? mem_1842 : _GEN_1846;
  assign _GEN_1848 = 11'h733 == _T_12323 ? mem_1843 : _GEN_1847;
  assign _GEN_1849 = 11'h734 == _T_12323 ? mem_1844 : _GEN_1848;
  assign _GEN_1850 = 11'h735 == _T_12323 ? mem_1845 : _GEN_1849;
  assign _GEN_1851 = 11'h736 == _T_12323 ? mem_1846 : _GEN_1850;
  assign _GEN_1852 = 11'h737 == _T_12323 ? mem_1847 : _GEN_1851;
  assign _GEN_1853 = 11'h738 == _T_12323 ? mem_1848 : _GEN_1852;
  assign _GEN_1854 = 11'h739 == _T_12323 ? mem_1849 : _GEN_1853;
  assign _GEN_1855 = 11'h73a == _T_12323 ? mem_1850 : _GEN_1854;
  assign _GEN_1856 = 11'h73b == _T_12323 ? mem_1851 : _GEN_1855;
  assign _GEN_1857 = 11'h73c == _T_12323 ? mem_1852 : _GEN_1856;
  assign _GEN_1858 = 11'h73d == _T_12323 ? mem_1853 : _GEN_1857;
  assign _GEN_1859 = 11'h73e == _T_12323 ? mem_1854 : _GEN_1858;
  assign _GEN_1860 = 11'h73f == _T_12323 ? mem_1855 : _GEN_1859;
  assign _GEN_1861 = 11'h740 == _T_12323 ? mem_1856 : _GEN_1860;
  assign _GEN_1862 = 11'h741 == _T_12323 ? mem_1857 : _GEN_1861;
  assign _GEN_1863 = 11'h742 == _T_12323 ? mem_1858 : _GEN_1862;
  assign _GEN_1864 = 11'h743 == _T_12323 ? mem_1859 : _GEN_1863;
  assign _GEN_1865 = 11'h744 == _T_12323 ? mem_1860 : _GEN_1864;
  assign _GEN_1866 = 11'h745 == _T_12323 ? mem_1861 : _GEN_1865;
  assign _GEN_1867 = 11'h746 == _T_12323 ? mem_1862 : _GEN_1866;
  assign _GEN_1868 = 11'h747 == _T_12323 ? mem_1863 : _GEN_1867;
  assign _GEN_1869 = 11'h748 == _T_12323 ? mem_1864 : _GEN_1868;
  assign _GEN_1870 = 11'h749 == _T_12323 ? mem_1865 : _GEN_1869;
  assign _GEN_1871 = 11'h74a == _T_12323 ? mem_1866 : _GEN_1870;
  assign _GEN_1872 = 11'h74b == _T_12323 ? mem_1867 : _GEN_1871;
  assign _GEN_1873 = 11'h74c == _T_12323 ? mem_1868 : _GEN_1872;
  assign _GEN_1874 = 11'h74d == _T_12323 ? mem_1869 : _GEN_1873;
  assign _GEN_1875 = 11'h74e == _T_12323 ? mem_1870 : _GEN_1874;
  assign _GEN_1876 = 11'h74f == _T_12323 ? mem_1871 : _GEN_1875;
  assign _GEN_1877 = 11'h750 == _T_12323 ? mem_1872 : _GEN_1876;
  assign _GEN_1878 = 11'h751 == _T_12323 ? mem_1873 : _GEN_1877;
  assign _GEN_1879 = 11'h752 == _T_12323 ? mem_1874 : _GEN_1878;
  assign _GEN_1880 = 11'h753 == _T_12323 ? mem_1875 : _GEN_1879;
  assign _GEN_1881 = 11'h754 == _T_12323 ? mem_1876 : _GEN_1880;
  assign _GEN_1882 = 11'h755 == _T_12323 ? mem_1877 : _GEN_1881;
  assign _GEN_1883 = 11'h756 == _T_12323 ? mem_1878 : _GEN_1882;
  assign _GEN_1884 = 11'h757 == _T_12323 ? mem_1879 : _GEN_1883;
  assign _GEN_1885 = 11'h758 == _T_12323 ? mem_1880 : _GEN_1884;
  assign _GEN_1886 = 11'h759 == _T_12323 ? mem_1881 : _GEN_1885;
  assign _GEN_1887 = 11'h75a == _T_12323 ? mem_1882 : _GEN_1886;
  assign _GEN_1888 = 11'h75b == _T_12323 ? mem_1883 : _GEN_1887;
  assign _GEN_1889 = 11'h75c == _T_12323 ? mem_1884 : _GEN_1888;
  assign _GEN_1890 = 11'h75d == _T_12323 ? mem_1885 : _GEN_1889;
  assign _GEN_1891 = 11'h75e == _T_12323 ? mem_1886 : _GEN_1890;
  assign _GEN_1892 = 11'h75f == _T_12323 ? mem_1887 : _GEN_1891;
  assign _GEN_1893 = 11'h760 == _T_12323 ? mem_1888 : _GEN_1892;
  assign _GEN_1894 = 11'h761 == _T_12323 ? mem_1889 : _GEN_1893;
  assign _GEN_1895 = 11'h762 == _T_12323 ? mem_1890 : _GEN_1894;
  assign _GEN_1896 = 11'h763 == _T_12323 ? mem_1891 : _GEN_1895;
  assign _GEN_1897 = 11'h764 == _T_12323 ? mem_1892 : _GEN_1896;
  assign _GEN_1898 = 11'h765 == _T_12323 ? mem_1893 : _GEN_1897;
  assign _GEN_1899 = 11'h766 == _T_12323 ? mem_1894 : _GEN_1898;
  assign _GEN_1900 = 11'h767 == _T_12323 ? mem_1895 : _GEN_1899;
  assign _GEN_1901 = 11'h768 == _T_12323 ? mem_1896 : _GEN_1900;
  assign _GEN_1902 = 11'h769 == _T_12323 ? mem_1897 : _GEN_1901;
  assign _GEN_1903 = 11'h76a == _T_12323 ? mem_1898 : _GEN_1902;
  assign _GEN_1904 = 11'h76b == _T_12323 ? mem_1899 : _GEN_1903;
  assign _GEN_1905 = 11'h76c == _T_12323 ? mem_1900 : _GEN_1904;
  assign _GEN_1906 = 11'h76d == _T_12323 ? mem_1901 : _GEN_1905;
  assign _GEN_1907 = 11'h76e == _T_12323 ? mem_1902 : _GEN_1906;
  assign _GEN_1908 = 11'h76f == _T_12323 ? mem_1903 : _GEN_1907;
  assign _GEN_1909 = 11'h770 == _T_12323 ? mem_1904 : _GEN_1908;
  assign _GEN_1910 = 11'h771 == _T_12323 ? mem_1905 : _GEN_1909;
  assign _GEN_1911 = 11'h772 == _T_12323 ? mem_1906 : _GEN_1910;
  assign _GEN_1912 = 11'h773 == _T_12323 ? mem_1907 : _GEN_1911;
  assign _GEN_1913 = 11'h774 == _T_12323 ? mem_1908 : _GEN_1912;
  assign _GEN_1914 = 11'h775 == _T_12323 ? mem_1909 : _GEN_1913;
  assign _GEN_1915 = 11'h776 == _T_12323 ? mem_1910 : _GEN_1914;
  assign _GEN_1916 = 11'h777 == _T_12323 ? mem_1911 : _GEN_1915;
  assign _GEN_1917 = 11'h778 == _T_12323 ? mem_1912 : _GEN_1916;
  assign _GEN_1918 = 11'h779 == _T_12323 ? mem_1913 : _GEN_1917;
  assign _GEN_1919 = 11'h77a == _T_12323 ? mem_1914 : _GEN_1918;
  assign _GEN_1920 = 11'h77b == _T_12323 ? mem_1915 : _GEN_1919;
  assign _GEN_1921 = 11'h77c == _T_12323 ? mem_1916 : _GEN_1920;
  assign _GEN_1922 = 11'h77d == _T_12323 ? mem_1917 : _GEN_1921;
  assign _GEN_1923 = 11'h77e == _T_12323 ? mem_1918 : _GEN_1922;
  assign _GEN_1924 = 11'h77f == _T_12323 ? mem_1919 : _GEN_1923;
  assign _GEN_1925 = 11'h780 == _T_12323 ? mem_1920 : _GEN_1924;
  assign _GEN_1926 = 11'h781 == _T_12323 ? mem_1921 : _GEN_1925;
  assign _GEN_1927 = 11'h782 == _T_12323 ? mem_1922 : _GEN_1926;
  assign _GEN_1928 = 11'h783 == _T_12323 ? mem_1923 : _GEN_1927;
  assign _GEN_1929 = 11'h784 == _T_12323 ? mem_1924 : _GEN_1928;
  assign _GEN_1930 = 11'h785 == _T_12323 ? mem_1925 : _GEN_1929;
  assign _GEN_1931 = 11'h786 == _T_12323 ? mem_1926 : _GEN_1930;
  assign _GEN_1932 = 11'h787 == _T_12323 ? mem_1927 : _GEN_1931;
  assign _GEN_1933 = 11'h788 == _T_12323 ? mem_1928 : _GEN_1932;
  assign _GEN_1934 = 11'h789 == _T_12323 ? mem_1929 : _GEN_1933;
  assign _GEN_1935 = 11'h78a == _T_12323 ? mem_1930 : _GEN_1934;
  assign _GEN_1936 = 11'h78b == _T_12323 ? mem_1931 : _GEN_1935;
  assign _GEN_1937 = 11'h78c == _T_12323 ? mem_1932 : _GEN_1936;
  assign _GEN_1938 = 11'h78d == _T_12323 ? mem_1933 : _GEN_1937;
  assign _GEN_1939 = 11'h78e == _T_12323 ? mem_1934 : _GEN_1938;
  assign _GEN_1940 = 11'h78f == _T_12323 ? mem_1935 : _GEN_1939;
  assign _GEN_1941 = 11'h790 == _T_12323 ? mem_1936 : _GEN_1940;
  assign _GEN_1942 = 11'h791 == _T_12323 ? mem_1937 : _GEN_1941;
  assign _GEN_1943 = 11'h792 == _T_12323 ? mem_1938 : _GEN_1942;
  assign _GEN_1944 = 11'h793 == _T_12323 ? mem_1939 : _GEN_1943;
  assign _GEN_1945 = 11'h794 == _T_12323 ? mem_1940 : _GEN_1944;
  assign _GEN_1946 = 11'h795 == _T_12323 ? mem_1941 : _GEN_1945;
  assign _GEN_1947 = 11'h796 == _T_12323 ? mem_1942 : _GEN_1946;
  assign _GEN_1948 = 11'h797 == _T_12323 ? mem_1943 : _GEN_1947;
  assign _GEN_1949 = 11'h798 == _T_12323 ? mem_1944 : _GEN_1948;
  assign _GEN_1950 = 11'h799 == _T_12323 ? mem_1945 : _GEN_1949;
  assign _GEN_1951 = 11'h79a == _T_12323 ? mem_1946 : _GEN_1950;
  assign _GEN_1952 = 11'h79b == _T_12323 ? mem_1947 : _GEN_1951;
  assign _GEN_1953 = 11'h79c == _T_12323 ? mem_1948 : _GEN_1952;
  assign _GEN_1954 = 11'h79d == _T_12323 ? mem_1949 : _GEN_1953;
  assign _GEN_1955 = 11'h79e == _T_12323 ? mem_1950 : _GEN_1954;
  assign _GEN_1956 = 11'h79f == _T_12323 ? mem_1951 : _GEN_1955;
  assign _GEN_1957 = 11'h7a0 == _T_12323 ? mem_1952 : _GEN_1956;
  assign _GEN_1958 = 11'h7a1 == _T_12323 ? mem_1953 : _GEN_1957;
  assign _GEN_1959 = 11'h7a2 == _T_12323 ? mem_1954 : _GEN_1958;
  assign _GEN_1960 = 11'h7a3 == _T_12323 ? mem_1955 : _GEN_1959;
  assign _GEN_1961 = 11'h7a4 == _T_12323 ? mem_1956 : _GEN_1960;
  assign _GEN_1962 = 11'h7a5 == _T_12323 ? mem_1957 : _GEN_1961;
  assign _GEN_1963 = 11'h7a6 == _T_12323 ? mem_1958 : _GEN_1962;
  assign _GEN_1964 = 11'h7a7 == _T_12323 ? mem_1959 : _GEN_1963;
  assign _GEN_1965 = 11'h7a8 == _T_12323 ? mem_1960 : _GEN_1964;
  assign _GEN_1966 = 11'h7a9 == _T_12323 ? mem_1961 : _GEN_1965;
  assign _GEN_1967 = 11'h7aa == _T_12323 ? mem_1962 : _GEN_1966;
  assign _GEN_1968 = 11'h7ab == _T_12323 ? mem_1963 : _GEN_1967;
  assign _GEN_1969 = 11'h7ac == _T_12323 ? mem_1964 : _GEN_1968;
  assign _GEN_1970 = 11'h7ad == _T_12323 ? mem_1965 : _GEN_1969;
  assign _GEN_1971 = 11'h7ae == _T_12323 ? mem_1966 : _GEN_1970;
  assign _GEN_1972 = 11'h7af == _T_12323 ? mem_1967 : _GEN_1971;
  assign _GEN_1973 = 11'h7b0 == _T_12323 ? mem_1968 : _GEN_1972;
  assign _GEN_1974 = 11'h7b1 == _T_12323 ? mem_1969 : _GEN_1973;
  assign _GEN_1975 = 11'h7b2 == _T_12323 ? mem_1970 : _GEN_1974;
  assign _GEN_1976 = 11'h7b3 == _T_12323 ? mem_1971 : _GEN_1975;
  assign _GEN_1977 = 11'h7b4 == _T_12323 ? mem_1972 : _GEN_1976;
  assign _GEN_1978 = 11'h7b5 == _T_12323 ? mem_1973 : _GEN_1977;
  assign _GEN_1979 = 11'h7b6 == _T_12323 ? mem_1974 : _GEN_1978;
  assign _GEN_1980 = 11'h7b7 == _T_12323 ? mem_1975 : _GEN_1979;
  assign _GEN_1981 = 11'h7b8 == _T_12323 ? mem_1976 : _GEN_1980;
  assign _GEN_1982 = 11'h7b9 == _T_12323 ? mem_1977 : _GEN_1981;
  assign _GEN_1983 = 11'h7ba == _T_12323 ? mem_1978 : _GEN_1982;
  assign _GEN_1984 = 11'h7bb == _T_12323 ? mem_1979 : _GEN_1983;
  assign _GEN_1985 = 11'h7bc == _T_12323 ? mem_1980 : _GEN_1984;
  assign _GEN_1986 = 11'h7bd == _T_12323 ? mem_1981 : _GEN_1985;
  assign _GEN_1987 = 11'h7be == _T_12323 ? mem_1982 : _GEN_1986;
  assign _GEN_1988 = 11'h7bf == _T_12323 ? mem_1983 : _GEN_1987;
  assign _GEN_1989 = 11'h7c0 == _T_12323 ? mem_1984 : _GEN_1988;
  assign _GEN_1990 = 11'h7c1 == _T_12323 ? mem_1985 : _GEN_1989;
  assign _GEN_1991 = 11'h7c2 == _T_12323 ? mem_1986 : _GEN_1990;
  assign _GEN_1992 = 11'h7c3 == _T_12323 ? mem_1987 : _GEN_1991;
  assign _GEN_1993 = 11'h7c4 == _T_12323 ? mem_1988 : _GEN_1992;
  assign _GEN_1994 = 11'h7c5 == _T_12323 ? mem_1989 : _GEN_1993;
  assign _GEN_1995 = 11'h7c6 == _T_12323 ? mem_1990 : _GEN_1994;
  assign _GEN_1996 = 11'h7c7 == _T_12323 ? mem_1991 : _GEN_1995;
  assign _GEN_1997 = 11'h7c8 == _T_12323 ? mem_1992 : _GEN_1996;
  assign _GEN_1998 = 11'h7c9 == _T_12323 ? mem_1993 : _GEN_1997;
  assign _GEN_1999 = 11'h7ca == _T_12323 ? mem_1994 : _GEN_1998;
  assign _GEN_2000 = 11'h7cb == _T_12323 ? mem_1995 : _GEN_1999;
  assign _GEN_2001 = 11'h7cc == _T_12323 ? mem_1996 : _GEN_2000;
  assign _GEN_2002 = 11'h7cd == _T_12323 ? mem_1997 : _GEN_2001;
  assign _GEN_2003 = 11'h7ce == _T_12323 ? mem_1998 : _GEN_2002;
  assign _GEN_2004 = 11'h7cf == _T_12323 ? mem_1999 : _GEN_2003;
  assign _GEN_2005 = 11'h7d0 == _T_12323 ? mem_2000 : _GEN_2004;
  assign _GEN_2006 = 11'h7d1 == _T_12323 ? mem_2001 : _GEN_2005;
  assign _GEN_2007 = 11'h7d2 == _T_12323 ? mem_2002 : _GEN_2006;
  assign _GEN_2008 = 11'h7d3 == _T_12323 ? mem_2003 : _GEN_2007;
  assign _GEN_2009 = 11'h7d4 == _T_12323 ? mem_2004 : _GEN_2008;
  assign _GEN_2010 = 11'h7d5 == _T_12323 ? mem_2005 : _GEN_2009;
  assign _GEN_2011 = 11'h7d6 == _T_12323 ? mem_2006 : _GEN_2010;
  assign _GEN_2012 = 11'h7d7 == _T_12323 ? mem_2007 : _GEN_2011;
  assign _GEN_2013 = 11'h7d8 == _T_12323 ? mem_2008 : _GEN_2012;
  assign _GEN_2014 = 11'h7d9 == _T_12323 ? mem_2009 : _GEN_2013;
  assign _GEN_2015 = 11'h7da == _T_12323 ? mem_2010 : _GEN_2014;
  assign _GEN_2016 = 11'h7db == _T_12323 ? mem_2011 : _GEN_2015;
  assign _GEN_2017 = 11'h7dc == _T_12323 ? mem_2012 : _GEN_2016;
  assign _GEN_2018 = 11'h7dd == _T_12323 ? mem_2013 : _GEN_2017;
  assign _GEN_2019 = 11'h7de == _T_12323 ? mem_2014 : _GEN_2018;
  assign _GEN_2020 = 11'h7df == _T_12323 ? mem_2015 : _GEN_2019;
  assign _GEN_2021 = 11'h7e0 == _T_12323 ? mem_2016 : _GEN_2020;
  assign _GEN_2022 = 11'h7e1 == _T_12323 ? mem_2017 : _GEN_2021;
  assign _GEN_2023 = 11'h7e2 == _T_12323 ? mem_2018 : _GEN_2022;
  assign _GEN_2024 = 11'h7e3 == _T_12323 ? mem_2019 : _GEN_2023;
  assign _GEN_2025 = 11'h7e4 == _T_12323 ? mem_2020 : _GEN_2024;
  assign _GEN_2026 = 11'h7e5 == _T_12323 ? mem_2021 : _GEN_2025;
  assign _GEN_2027 = 11'h7e6 == _T_12323 ? mem_2022 : _GEN_2026;
  assign _GEN_2028 = 11'h7e7 == _T_12323 ? mem_2023 : _GEN_2027;
  assign _GEN_2029 = 11'h7e8 == _T_12323 ? mem_2024 : _GEN_2028;
  assign _GEN_2030 = 11'h7e9 == _T_12323 ? mem_2025 : _GEN_2029;
  assign _GEN_2031 = 11'h7ea == _T_12323 ? mem_2026 : _GEN_2030;
  assign _GEN_2032 = 11'h7eb == _T_12323 ? mem_2027 : _GEN_2031;
  assign _GEN_2033 = 11'h7ec == _T_12323 ? mem_2028 : _GEN_2032;
  assign _GEN_2034 = 11'h7ed == _T_12323 ? mem_2029 : _GEN_2033;
  assign _GEN_2035 = 11'h7ee == _T_12323 ? mem_2030 : _GEN_2034;
  assign _GEN_2036 = 11'h7ef == _T_12323 ? mem_2031 : _GEN_2035;
  assign _GEN_2037 = 11'h7f0 == _T_12323 ? mem_2032 : _GEN_2036;
  assign _GEN_2038 = 11'h7f1 == _T_12323 ? mem_2033 : _GEN_2037;
  assign _GEN_2039 = 11'h7f2 == _T_12323 ? mem_2034 : _GEN_2038;
  assign _GEN_2040 = 11'h7f3 == _T_12323 ? mem_2035 : _GEN_2039;
  assign _GEN_2041 = 11'h7f4 == _T_12323 ? mem_2036 : _GEN_2040;
  assign _GEN_2042 = 11'h7f5 == _T_12323 ? mem_2037 : _GEN_2041;
  assign _GEN_2043 = 11'h7f6 == _T_12323 ? mem_2038 : _GEN_2042;
  assign _GEN_2044 = 11'h7f7 == _T_12323 ? mem_2039 : _GEN_2043;
  assign _GEN_2045 = 11'h7f8 == _T_12323 ? mem_2040 : _GEN_2044;
  assign _GEN_2046 = 11'h7f9 == _T_12323 ? mem_2041 : _GEN_2045;
  assign _GEN_2047 = 11'h7fa == _T_12323 ? mem_2042 : _GEN_2046;
  assign _GEN_2048 = 11'h7fb == _T_12323 ? mem_2043 : _GEN_2047;
  assign _GEN_2049 = 11'h7fc == _T_12323 ? mem_2044 : _GEN_2048;
  assign _GEN_2050 = 11'h7fd == _T_12323 ? mem_2045 : _GEN_2049;
  assign _GEN_2051 = 11'h7fe == _T_12323 ? mem_2046 : _GEN_2050;
  assign _GEN_2052 = 11'h7ff == _T_12323 ? mem_2047 : _GEN_2051;
  assign _T_12324 = _GEN_0[7:0];
  assign _GEN_2053 = _T_12316 ? _T_12319 : _T_12324;
  assign _T_12325 = wen[1];
  assign _T_12328 = wdata[15:8];
  assign _T_12333 = _GEN_1[15:8];
  assign _GEN_4101 = _T_12325 ? _T_12328 : _T_12333;
  assign _T_12334 = wen[2];
  assign _T_12337 = wdata[23:16];
  assign _T_12342 = _GEN_2[23:16];
  assign _GEN_6149 = _T_12334 ? _T_12337 : _T_12342;
  assign _T_12343 = wen[3];
  assign _T_12346 = wdata[31:24];
  assign _T_12351 = _GEN_3[31:24];
  assign _GEN_8197 = _T_12343 ? _T_12346 : _T_12351;
  assign _T_12356 = {toWrite_1,toWrite_0};
  assign _T_12357 = {toWrite_2,_T_12356};
  assign _T_12358 = {toWrite_3,_T_12357};
  assign _GEN_8198 = 11'h0 == _T_12323 ? _GEN_4 : mem_0;
  assign _GEN_8199 = 11'h1 == _T_12323 ? _GEN_4 : mem_1;
  assign _GEN_8200 = 11'h2 == _T_12323 ? _GEN_4 : mem_2;
  assign _GEN_8201 = 11'h3 == _T_12323 ? _GEN_4 : mem_3;
  assign _GEN_8202 = 11'h4 == _T_12323 ? _GEN_4 : mem_4;
  assign _GEN_8203 = 11'h5 == _T_12323 ? _GEN_4 : mem_5;
  assign _GEN_8204 = 11'h6 == _T_12323 ? _GEN_4 : mem_6;
  assign _GEN_8205 = 11'h7 == _T_12323 ? _GEN_4 : mem_7;
  assign _GEN_8206 = 11'h8 == _T_12323 ? _GEN_4 : mem_8;
  assign _GEN_8207 = 11'h9 == _T_12323 ? _GEN_4 : mem_9;
  assign _GEN_8208 = 11'ha == _T_12323 ? _GEN_4 : mem_10;
  assign _GEN_8209 = 11'hb == _T_12323 ? _GEN_4 : mem_11;
  assign _GEN_8210 = 11'hc == _T_12323 ? _GEN_4 : mem_12;
  assign _GEN_8211 = 11'hd == _T_12323 ? _GEN_4 : mem_13;
  assign _GEN_8212 = 11'he == _T_12323 ? _GEN_4 : mem_14;
  assign _GEN_8213 = 11'hf == _T_12323 ? _GEN_4 : mem_15;
  assign _GEN_8214 = 11'h10 == _T_12323 ? _GEN_4 : mem_16;
  assign _GEN_8215 = 11'h11 == _T_12323 ? _GEN_4 : mem_17;
  assign _GEN_8216 = 11'h12 == _T_12323 ? _GEN_4 : mem_18;
  assign _GEN_8217 = 11'h13 == _T_12323 ? _GEN_4 : mem_19;
  assign _GEN_8218 = 11'h14 == _T_12323 ? _GEN_4 : mem_20;
  assign _GEN_8219 = 11'h15 == _T_12323 ? _GEN_4 : mem_21;
  assign _GEN_8220 = 11'h16 == _T_12323 ? _GEN_4 : mem_22;
  assign _GEN_8221 = 11'h17 == _T_12323 ? _GEN_4 : mem_23;
  assign _GEN_8222 = 11'h18 == _T_12323 ? _GEN_4 : mem_24;
  assign _GEN_8223 = 11'h19 == _T_12323 ? _GEN_4 : mem_25;
  assign _GEN_8224 = 11'h1a == _T_12323 ? _GEN_4 : mem_26;
  assign _GEN_8225 = 11'h1b == _T_12323 ? _GEN_4 : mem_27;
  assign _GEN_8226 = 11'h1c == _T_12323 ? _GEN_4 : mem_28;
  assign _GEN_8227 = 11'h1d == _T_12323 ? _GEN_4 : mem_29;
  assign _GEN_8228 = 11'h1e == _T_12323 ? _GEN_4 : mem_30;
  assign _GEN_8229 = 11'h1f == _T_12323 ? _GEN_4 : mem_31;
  assign _GEN_8230 = 11'h20 == _T_12323 ? _GEN_4 : mem_32;
  assign _GEN_8231 = 11'h21 == _T_12323 ? _GEN_4 : mem_33;
  assign _GEN_8232 = 11'h22 == _T_12323 ? _GEN_4 : mem_34;
  assign _GEN_8233 = 11'h23 == _T_12323 ? _GEN_4 : mem_35;
  assign _GEN_8234 = 11'h24 == _T_12323 ? _GEN_4 : mem_36;
  assign _GEN_8235 = 11'h25 == _T_12323 ? _GEN_4 : mem_37;
  assign _GEN_8236 = 11'h26 == _T_12323 ? _GEN_4 : mem_38;
  assign _GEN_8237 = 11'h27 == _T_12323 ? _GEN_4 : mem_39;
  assign _GEN_8238 = 11'h28 == _T_12323 ? _GEN_4 : mem_40;
  assign _GEN_8239 = 11'h29 == _T_12323 ? _GEN_4 : mem_41;
  assign _GEN_8240 = 11'h2a == _T_12323 ? _GEN_4 : mem_42;
  assign _GEN_8241 = 11'h2b == _T_12323 ? _GEN_4 : mem_43;
  assign _GEN_8242 = 11'h2c == _T_12323 ? _GEN_4 : mem_44;
  assign _GEN_8243 = 11'h2d == _T_12323 ? _GEN_4 : mem_45;
  assign _GEN_8244 = 11'h2e == _T_12323 ? _GEN_4 : mem_46;
  assign _GEN_8245 = 11'h2f == _T_12323 ? _GEN_4 : mem_47;
  assign _GEN_8246 = 11'h30 == _T_12323 ? _GEN_4 : mem_48;
  assign _GEN_8247 = 11'h31 == _T_12323 ? _GEN_4 : mem_49;
  assign _GEN_8248 = 11'h32 == _T_12323 ? _GEN_4 : mem_50;
  assign _GEN_8249 = 11'h33 == _T_12323 ? _GEN_4 : mem_51;
  assign _GEN_8250 = 11'h34 == _T_12323 ? _GEN_4 : mem_52;
  assign _GEN_8251 = 11'h35 == _T_12323 ? _GEN_4 : mem_53;
  assign _GEN_8252 = 11'h36 == _T_12323 ? _GEN_4 : mem_54;
  assign _GEN_8253 = 11'h37 == _T_12323 ? _GEN_4 : mem_55;
  assign _GEN_8254 = 11'h38 == _T_12323 ? _GEN_4 : mem_56;
  assign _GEN_8255 = 11'h39 == _T_12323 ? _GEN_4 : mem_57;
  assign _GEN_8256 = 11'h3a == _T_12323 ? _GEN_4 : mem_58;
  assign _GEN_8257 = 11'h3b == _T_12323 ? _GEN_4 : mem_59;
  assign _GEN_8258 = 11'h3c == _T_12323 ? _GEN_4 : mem_60;
  assign _GEN_8259 = 11'h3d == _T_12323 ? _GEN_4 : mem_61;
  assign _GEN_8260 = 11'h3e == _T_12323 ? _GEN_4 : mem_62;
  assign _GEN_8261 = 11'h3f == _T_12323 ? _GEN_4 : mem_63;
  assign _GEN_8262 = 11'h40 == _T_12323 ? _GEN_4 : mem_64;
  assign _GEN_8263 = 11'h41 == _T_12323 ? _GEN_4 : mem_65;
  assign _GEN_8264 = 11'h42 == _T_12323 ? _GEN_4 : mem_66;
  assign _GEN_8265 = 11'h43 == _T_12323 ? _GEN_4 : mem_67;
  assign _GEN_8266 = 11'h44 == _T_12323 ? _GEN_4 : mem_68;
  assign _GEN_8267 = 11'h45 == _T_12323 ? _GEN_4 : mem_69;
  assign _GEN_8268 = 11'h46 == _T_12323 ? _GEN_4 : mem_70;
  assign _GEN_8269 = 11'h47 == _T_12323 ? _GEN_4 : mem_71;
  assign _GEN_8270 = 11'h48 == _T_12323 ? _GEN_4 : mem_72;
  assign _GEN_8271 = 11'h49 == _T_12323 ? _GEN_4 : mem_73;
  assign _GEN_8272 = 11'h4a == _T_12323 ? _GEN_4 : mem_74;
  assign _GEN_8273 = 11'h4b == _T_12323 ? _GEN_4 : mem_75;
  assign _GEN_8274 = 11'h4c == _T_12323 ? _GEN_4 : mem_76;
  assign _GEN_8275 = 11'h4d == _T_12323 ? _GEN_4 : mem_77;
  assign _GEN_8276 = 11'h4e == _T_12323 ? _GEN_4 : mem_78;
  assign _GEN_8277 = 11'h4f == _T_12323 ? _GEN_4 : mem_79;
  assign _GEN_8278 = 11'h50 == _T_12323 ? _GEN_4 : mem_80;
  assign _GEN_8279 = 11'h51 == _T_12323 ? _GEN_4 : mem_81;
  assign _GEN_8280 = 11'h52 == _T_12323 ? _GEN_4 : mem_82;
  assign _GEN_8281 = 11'h53 == _T_12323 ? _GEN_4 : mem_83;
  assign _GEN_8282 = 11'h54 == _T_12323 ? _GEN_4 : mem_84;
  assign _GEN_8283 = 11'h55 == _T_12323 ? _GEN_4 : mem_85;
  assign _GEN_8284 = 11'h56 == _T_12323 ? _GEN_4 : mem_86;
  assign _GEN_8285 = 11'h57 == _T_12323 ? _GEN_4 : mem_87;
  assign _GEN_8286 = 11'h58 == _T_12323 ? _GEN_4 : mem_88;
  assign _GEN_8287 = 11'h59 == _T_12323 ? _GEN_4 : mem_89;
  assign _GEN_8288 = 11'h5a == _T_12323 ? _GEN_4 : mem_90;
  assign _GEN_8289 = 11'h5b == _T_12323 ? _GEN_4 : mem_91;
  assign _GEN_8290 = 11'h5c == _T_12323 ? _GEN_4 : mem_92;
  assign _GEN_8291 = 11'h5d == _T_12323 ? _GEN_4 : mem_93;
  assign _GEN_8292 = 11'h5e == _T_12323 ? _GEN_4 : mem_94;
  assign _GEN_8293 = 11'h5f == _T_12323 ? _GEN_4 : mem_95;
  assign _GEN_8294 = 11'h60 == _T_12323 ? _GEN_4 : mem_96;
  assign _GEN_8295 = 11'h61 == _T_12323 ? _GEN_4 : mem_97;
  assign _GEN_8296 = 11'h62 == _T_12323 ? _GEN_4 : mem_98;
  assign _GEN_8297 = 11'h63 == _T_12323 ? _GEN_4 : mem_99;
  assign _GEN_8298 = 11'h64 == _T_12323 ? _GEN_4 : mem_100;
  assign _GEN_8299 = 11'h65 == _T_12323 ? _GEN_4 : mem_101;
  assign _GEN_8300 = 11'h66 == _T_12323 ? _GEN_4 : mem_102;
  assign _GEN_8301 = 11'h67 == _T_12323 ? _GEN_4 : mem_103;
  assign _GEN_8302 = 11'h68 == _T_12323 ? _GEN_4 : mem_104;
  assign _GEN_8303 = 11'h69 == _T_12323 ? _GEN_4 : mem_105;
  assign _GEN_8304 = 11'h6a == _T_12323 ? _GEN_4 : mem_106;
  assign _GEN_8305 = 11'h6b == _T_12323 ? _GEN_4 : mem_107;
  assign _GEN_8306 = 11'h6c == _T_12323 ? _GEN_4 : mem_108;
  assign _GEN_8307 = 11'h6d == _T_12323 ? _GEN_4 : mem_109;
  assign _GEN_8308 = 11'h6e == _T_12323 ? _GEN_4 : mem_110;
  assign _GEN_8309 = 11'h6f == _T_12323 ? _GEN_4 : mem_111;
  assign _GEN_8310 = 11'h70 == _T_12323 ? _GEN_4 : mem_112;
  assign _GEN_8311 = 11'h71 == _T_12323 ? _GEN_4 : mem_113;
  assign _GEN_8312 = 11'h72 == _T_12323 ? _GEN_4 : mem_114;
  assign _GEN_8313 = 11'h73 == _T_12323 ? _GEN_4 : mem_115;
  assign _GEN_8314 = 11'h74 == _T_12323 ? _GEN_4 : mem_116;
  assign _GEN_8315 = 11'h75 == _T_12323 ? _GEN_4 : mem_117;
  assign _GEN_8316 = 11'h76 == _T_12323 ? _GEN_4 : mem_118;
  assign _GEN_8317 = 11'h77 == _T_12323 ? _GEN_4 : mem_119;
  assign _GEN_8318 = 11'h78 == _T_12323 ? _GEN_4 : mem_120;
  assign _GEN_8319 = 11'h79 == _T_12323 ? _GEN_4 : mem_121;
  assign _GEN_8320 = 11'h7a == _T_12323 ? _GEN_4 : mem_122;
  assign _GEN_8321 = 11'h7b == _T_12323 ? _GEN_4 : mem_123;
  assign _GEN_8322 = 11'h7c == _T_12323 ? _GEN_4 : mem_124;
  assign _GEN_8323 = 11'h7d == _T_12323 ? _GEN_4 : mem_125;
  assign _GEN_8324 = 11'h7e == _T_12323 ? _GEN_4 : mem_126;
  assign _GEN_8325 = 11'h7f == _T_12323 ? _GEN_4 : mem_127;
  assign _GEN_8326 = 11'h80 == _T_12323 ? _GEN_4 : mem_128;
  assign _GEN_8327 = 11'h81 == _T_12323 ? _GEN_4 : mem_129;
  assign _GEN_8328 = 11'h82 == _T_12323 ? _GEN_4 : mem_130;
  assign _GEN_8329 = 11'h83 == _T_12323 ? _GEN_4 : mem_131;
  assign _GEN_8330 = 11'h84 == _T_12323 ? _GEN_4 : mem_132;
  assign _GEN_8331 = 11'h85 == _T_12323 ? _GEN_4 : mem_133;
  assign _GEN_8332 = 11'h86 == _T_12323 ? _GEN_4 : mem_134;
  assign _GEN_8333 = 11'h87 == _T_12323 ? _GEN_4 : mem_135;
  assign _GEN_8334 = 11'h88 == _T_12323 ? _GEN_4 : mem_136;
  assign _GEN_8335 = 11'h89 == _T_12323 ? _GEN_4 : mem_137;
  assign _GEN_8336 = 11'h8a == _T_12323 ? _GEN_4 : mem_138;
  assign _GEN_8337 = 11'h8b == _T_12323 ? _GEN_4 : mem_139;
  assign _GEN_8338 = 11'h8c == _T_12323 ? _GEN_4 : mem_140;
  assign _GEN_8339 = 11'h8d == _T_12323 ? _GEN_4 : mem_141;
  assign _GEN_8340 = 11'h8e == _T_12323 ? _GEN_4 : mem_142;
  assign _GEN_8341 = 11'h8f == _T_12323 ? _GEN_4 : mem_143;
  assign _GEN_8342 = 11'h90 == _T_12323 ? _GEN_4 : mem_144;
  assign _GEN_8343 = 11'h91 == _T_12323 ? _GEN_4 : mem_145;
  assign _GEN_8344 = 11'h92 == _T_12323 ? _GEN_4 : mem_146;
  assign _GEN_8345 = 11'h93 == _T_12323 ? _GEN_4 : mem_147;
  assign _GEN_8346 = 11'h94 == _T_12323 ? _GEN_4 : mem_148;
  assign _GEN_8347 = 11'h95 == _T_12323 ? _GEN_4 : mem_149;
  assign _GEN_8348 = 11'h96 == _T_12323 ? _GEN_4 : mem_150;
  assign _GEN_8349 = 11'h97 == _T_12323 ? _GEN_4 : mem_151;
  assign _GEN_8350 = 11'h98 == _T_12323 ? _GEN_4 : mem_152;
  assign _GEN_8351 = 11'h99 == _T_12323 ? _GEN_4 : mem_153;
  assign _GEN_8352 = 11'h9a == _T_12323 ? _GEN_4 : mem_154;
  assign _GEN_8353 = 11'h9b == _T_12323 ? _GEN_4 : mem_155;
  assign _GEN_8354 = 11'h9c == _T_12323 ? _GEN_4 : mem_156;
  assign _GEN_8355 = 11'h9d == _T_12323 ? _GEN_4 : mem_157;
  assign _GEN_8356 = 11'h9e == _T_12323 ? _GEN_4 : mem_158;
  assign _GEN_8357 = 11'h9f == _T_12323 ? _GEN_4 : mem_159;
  assign _GEN_8358 = 11'ha0 == _T_12323 ? _GEN_4 : mem_160;
  assign _GEN_8359 = 11'ha1 == _T_12323 ? _GEN_4 : mem_161;
  assign _GEN_8360 = 11'ha2 == _T_12323 ? _GEN_4 : mem_162;
  assign _GEN_8361 = 11'ha3 == _T_12323 ? _GEN_4 : mem_163;
  assign _GEN_8362 = 11'ha4 == _T_12323 ? _GEN_4 : mem_164;
  assign _GEN_8363 = 11'ha5 == _T_12323 ? _GEN_4 : mem_165;
  assign _GEN_8364 = 11'ha6 == _T_12323 ? _GEN_4 : mem_166;
  assign _GEN_8365 = 11'ha7 == _T_12323 ? _GEN_4 : mem_167;
  assign _GEN_8366 = 11'ha8 == _T_12323 ? _GEN_4 : mem_168;
  assign _GEN_8367 = 11'ha9 == _T_12323 ? _GEN_4 : mem_169;
  assign _GEN_8368 = 11'haa == _T_12323 ? _GEN_4 : mem_170;
  assign _GEN_8369 = 11'hab == _T_12323 ? _GEN_4 : mem_171;
  assign _GEN_8370 = 11'hac == _T_12323 ? _GEN_4 : mem_172;
  assign _GEN_8371 = 11'had == _T_12323 ? _GEN_4 : mem_173;
  assign _GEN_8372 = 11'hae == _T_12323 ? _GEN_4 : mem_174;
  assign _GEN_8373 = 11'haf == _T_12323 ? _GEN_4 : mem_175;
  assign _GEN_8374 = 11'hb0 == _T_12323 ? _GEN_4 : mem_176;
  assign _GEN_8375 = 11'hb1 == _T_12323 ? _GEN_4 : mem_177;
  assign _GEN_8376 = 11'hb2 == _T_12323 ? _GEN_4 : mem_178;
  assign _GEN_8377 = 11'hb3 == _T_12323 ? _GEN_4 : mem_179;
  assign _GEN_8378 = 11'hb4 == _T_12323 ? _GEN_4 : mem_180;
  assign _GEN_8379 = 11'hb5 == _T_12323 ? _GEN_4 : mem_181;
  assign _GEN_8380 = 11'hb6 == _T_12323 ? _GEN_4 : mem_182;
  assign _GEN_8381 = 11'hb7 == _T_12323 ? _GEN_4 : mem_183;
  assign _GEN_8382 = 11'hb8 == _T_12323 ? _GEN_4 : mem_184;
  assign _GEN_8383 = 11'hb9 == _T_12323 ? _GEN_4 : mem_185;
  assign _GEN_8384 = 11'hba == _T_12323 ? _GEN_4 : mem_186;
  assign _GEN_8385 = 11'hbb == _T_12323 ? _GEN_4 : mem_187;
  assign _GEN_8386 = 11'hbc == _T_12323 ? _GEN_4 : mem_188;
  assign _GEN_8387 = 11'hbd == _T_12323 ? _GEN_4 : mem_189;
  assign _GEN_8388 = 11'hbe == _T_12323 ? _GEN_4 : mem_190;
  assign _GEN_8389 = 11'hbf == _T_12323 ? _GEN_4 : mem_191;
  assign _GEN_8390 = 11'hc0 == _T_12323 ? _GEN_4 : mem_192;
  assign _GEN_8391 = 11'hc1 == _T_12323 ? _GEN_4 : mem_193;
  assign _GEN_8392 = 11'hc2 == _T_12323 ? _GEN_4 : mem_194;
  assign _GEN_8393 = 11'hc3 == _T_12323 ? _GEN_4 : mem_195;
  assign _GEN_8394 = 11'hc4 == _T_12323 ? _GEN_4 : mem_196;
  assign _GEN_8395 = 11'hc5 == _T_12323 ? _GEN_4 : mem_197;
  assign _GEN_8396 = 11'hc6 == _T_12323 ? _GEN_4 : mem_198;
  assign _GEN_8397 = 11'hc7 == _T_12323 ? _GEN_4 : mem_199;
  assign _GEN_8398 = 11'hc8 == _T_12323 ? _GEN_4 : mem_200;
  assign _GEN_8399 = 11'hc9 == _T_12323 ? _GEN_4 : mem_201;
  assign _GEN_8400 = 11'hca == _T_12323 ? _GEN_4 : mem_202;
  assign _GEN_8401 = 11'hcb == _T_12323 ? _GEN_4 : mem_203;
  assign _GEN_8402 = 11'hcc == _T_12323 ? _GEN_4 : mem_204;
  assign _GEN_8403 = 11'hcd == _T_12323 ? _GEN_4 : mem_205;
  assign _GEN_8404 = 11'hce == _T_12323 ? _GEN_4 : mem_206;
  assign _GEN_8405 = 11'hcf == _T_12323 ? _GEN_4 : mem_207;
  assign _GEN_8406 = 11'hd0 == _T_12323 ? _GEN_4 : mem_208;
  assign _GEN_8407 = 11'hd1 == _T_12323 ? _GEN_4 : mem_209;
  assign _GEN_8408 = 11'hd2 == _T_12323 ? _GEN_4 : mem_210;
  assign _GEN_8409 = 11'hd3 == _T_12323 ? _GEN_4 : mem_211;
  assign _GEN_8410 = 11'hd4 == _T_12323 ? _GEN_4 : mem_212;
  assign _GEN_8411 = 11'hd5 == _T_12323 ? _GEN_4 : mem_213;
  assign _GEN_8412 = 11'hd6 == _T_12323 ? _GEN_4 : mem_214;
  assign _GEN_8413 = 11'hd7 == _T_12323 ? _GEN_4 : mem_215;
  assign _GEN_8414 = 11'hd8 == _T_12323 ? _GEN_4 : mem_216;
  assign _GEN_8415 = 11'hd9 == _T_12323 ? _GEN_4 : mem_217;
  assign _GEN_8416 = 11'hda == _T_12323 ? _GEN_4 : mem_218;
  assign _GEN_8417 = 11'hdb == _T_12323 ? _GEN_4 : mem_219;
  assign _GEN_8418 = 11'hdc == _T_12323 ? _GEN_4 : mem_220;
  assign _GEN_8419 = 11'hdd == _T_12323 ? _GEN_4 : mem_221;
  assign _GEN_8420 = 11'hde == _T_12323 ? _GEN_4 : mem_222;
  assign _GEN_8421 = 11'hdf == _T_12323 ? _GEN_4 : mem_223;
  assign _GEN_8422 = 11'he0 == _T_12323 ? _GEN_4 : mem_224;
  assign _GEN_8423 = 11'he1 == _T_12323 ? _GEN_4 : mem_225;
  assign _GEN_8424 = 11'he2 == _T_12323 ? _GEN_4 : mem_226;
  assign _GEN_8425 = 11'he3 == _T_12323 ? _GEN_4 : mem_227;
  assign _GEN_8426 = 11'he4 == _T_12323 ? _GEN_4 : mem_228;
  assign _GEN_8427 = 11'he5 == _T_12323 ? _GEN_4 : mem_229;
  assign _GEN_8428 = 11'he6 == _T_12323 ? _GEN_4 : mem_230;
  assign _GEN_8429 = 11'he7 == _T_12323 ? _GEN_4 : mem_231;
  assign _GEN_8430 = 11'he8 == _T_12323 ? _GEN_4 : mem_232;
  assign _GEN_8431 = 11'he9 == _T_12323 ? _GEN_4 : mem_233;
  assign _GEN_8432 = 11'hea == _T_12323 ? _GEN_4 : mem_234;
  assign _GEN_8433 = 11'heb == _T_12323 ? _GEN_4 : mem_235;
  assign _GEN_8434 = 11'hec == _T_12323 ? _GEN_4 : mem_236;
  assign _GEN_8435 = 11'hed == _T_12323 ? _GEN_4 : mem_237;
  assign _GEN_8436 = 11'hee == _T_12323 ? _GEN_4 : mem_238;
  assign _GEN_8437 = 11'hef == _T_12323 ? _GEN_4 : mem_239;
  assign _GEN_8438 = 11'hf0 == _T_12323 ? _GEN_4 : mem_240;
  assign _GEN_8439 = 11'hf1 == _T_12323 ? _GEN_4 : mem_241;
  assign _GEN_8440 = 11'hf2 == _T_12323 ? _GEN_4 : mem_242;
  assign _GEN_8441 = 11'hf3 == _T_12323 ? _GEN_4 : mem_243;
  assign _GEN_8442 = 11'hf4 == _T_12323 ? _GEN_4 : mem_244;
  assign _GEN_8443 = 11'hf5 == _T_12323 ? _GEN_4 : mem_245;
  assign _GEN_8444 = 11'hf6 == _T_12323 ? _GEN_4 : mem_246;
  assign _GEN_8445 = 11'hf7 == _T_12323 ? _GEN_4 : mem_247;
  assign _GEN_8446 = 11'hf8 == _T_12323 ? _GEN_4 : mem_248;
  assign _GEN_8447 = 11'hf9 == _T_12323 ? _GEN_4 : mem_249;
  assign _GEN_8448 = 11'hfa == _T_12323 ? _GEN_4 : mem_250;
  assign _GEN_8449 = 11'hfb == _T_12323 ? _GEN_4 : mem_251;
  assign _GEN_8450 = 11'hfc == _T_12323 ? _GEN_4 : mem_252;
  assign _GEN_8451 = 11'hfd == _T_12323 ? _GEN_4 : mem_253;
  assign _GEN_8452 = 11'hfe == _T_12323 ? _GEN_4 : mem_254;
  assign _GEN_8453 = 11'hff == _T_12323 ? _GEN_4 : mem_255;
  assign _GEN_8454 = 11'h100 == _T_12323 ? _GEN_4 : mem_256;
  assign _GEN_8455 = 11'h101 == _T_12323 ? _GEN_4 : mem_257;
  assign _GEN_8456 = 11'h102 == _T_12323 ? _GEN_4 : mem_258;
  assign _GEN_8457 = 11'h103 == _T_12323 ? _GEN_4 : mem_259;
  assign _GEN_8458 = 11'h104 == _T_12323 ? _GEN_4 : mem_260;
  assign _GEN_8459 = 11'h105 == _T_12323 ? _GEN_4 : mem_261;
  assign _GEN_8460 = 11'h106 == _T_12323 ? _GEN_4 : mem_262;
  assign _GEN_8461 = 11'h107 == _T_12323 ? _GEN_4 : mem_263;
  assign _GEN_8462 = 11'h108 == _T_12323 ? _GEN_4 : mem_264;
  assign _GEN_8463 = 11'h109 == _T_12323 ? _GEN_4 : mem_265;
  assign _GEN_8464 = 11'h10a == _T_12323 ? _GEN_4 : mem_266;
  assign _GEN_8465 = 11'h10b == _T_12323 ? _GEN_4 : mem_267;
  assign _GEN_8466 = 11'h10c == _T_12323 ? _GEN_4 : mem_268;
  assign _GEN_8467 = 11'h10d == _T_12323 ? _GEN_4 : mem_269;
  assign _GEN_8468 = 11'h10e == _T_12323 ? _GEN_4 : mem_270;
  assign _GEN_8469 = 11'h10f == _T_12323 ? _GEN_4 : mem_271;
  assign _GEN_8470 = 11'h110 == _T_12323 ? _GEN_4 : mem_272;
  assign _GEN_8471 = 11'h111 == _T_12323 ? _GEN_4 : mem_273;
  assign _GEN_8472 = 11'h112 == _T_12323 ? _GEN_4 : mem_274;
  assign _GEN_8473 = 11'h113 == _T_12323 ? _GEN_4 : mem_275;
  assign _GEN_8474 = 11'h114 == _T_12323 ? _GEN_4 : mem_276;
  assign _GEN_8475 = 11'h115 == _T_12323 ? _GEN_4 : mem_277;
  assign _GEN_8476 = 11'h116 == _T_12323 ? _GEN_4 : mem_278;
  assign _GEN_8477 = 11'h117 == _T_12323 ? _GEN_4 : mem_279;
  assign _GEN_8478 = 11'h118 == _T_12323 ? _GEN_4 : mem_280;
  assign _GEN_8479 = 11'h119 == _T_12323 ? _GEN_4 : mem_281;
  assign _GEN_8480 = 11'h11a == _T_12323 ? _GEN_4 : mem_282;
  assign _GEN_8481 = 11'h11b == _T_12323 ? _GEN_4 : mem_283;
  assign _GEN_8482 = 11'h11c == _T_12323 ? _GEN_4 : mem_284;
  assign _GEN_8483 = 11'h11d == _T_12323 ? _GEN_4 : mem_285;
  assign _GEN_8484 = 11'h11e == _T_12323 ? _GEN_4 : mem_286;
  assign _GEN_8485 = 11'h11f == _T_12323 ? _GEN_4 : mem_287;
  assign _GEN_8486 = 11'h120 == _T_12323 ? _GEN_4 : mem_288;
  assign _GEN_8487 = 11'h121 == _T_12323 ? _GEN_4 : mem_289;
  assign _GEN_8488 = 11'h122 == _T_12323 ? _GEN_4 : mem_290;
  assign _GEN_8489 = 11'h123 == _T_12323 ? _GEN_4 : mem_291;
  assign _GEN_8490 = 11'h124 == _T_12323 ? _GEN_4 : mem_292;
  assign _GEN_8491 = 11'h125 == _T_12323 ? _GEN_4 : mem_293;
  assign _GEN_8492 = 11'h126 == _T_12323 ? _GEN_4 : mem_294;
  assign _GEN_8493 = 11'h127 == _T_12323 ? _GEN_4 : mem_295;
  assign _GEN_8494 = 11'h128 == _T_12323 ? _GEN_4 : mem_296;
  assign _GEN_8495 = 11'h129 == _T_12323 ? _GEN_4 : mem_297;
  assign _GEN_8496 = 11'h12a == _T_12323 ? _GEN_4 : mem_298;
  assign _GEN_8497 = 11'h12b == _T_12323 ? _GEN_4 : mem_299;
  assign _GEN_8498 = 11'h12c == _T_12323 ? _GEN_4 : mem_300;
  assign _GEN_8499 = 11'h12d == _T_12323 ? _GEN_4 : mem_301;
  assign _GEN_8500 = 11'h12e == _T_12323 ? _GEN_4 : mem_302;
  assign _GEN_8501 = 11'h12f == _T_12323 ? _GEN_4 : mem_303;
  assign _GEN_8502 = 11'h130 == _T_12323 ? _GEN_4 : mem_304;
  assign _GEN_8503 = 11'h131 == _T_12323 ? _GEN_4 : mem_305;
  assign _GEN_8504 = 11'h132 == _T_12323 ? _GEN_4 : mem_306;
  assign _GEN_8505 = 11'h133 == _T_12323 ? _GEN_4 : mem_307;
  assign _GEN_8506 = 11'h134 == _T_12323 ? _GEN_4 : mem_308;
  assign _GEN_8507 = 11'h135 == _T_12323 ? _GEN_4 : mem_309;
  assign _GEN_8508 = 11'h136 == _T_12323 ? _GEN_4 : mem_310;
  assign _GEN_8509 = 11'h137 == _T_12323 ? _GEN_4 : mem_311;
  assign _GEN_8510 = 11'h138 == _T_12323 ? _GEN_4 : mem_312;
  assign _GEN_8511 = 11'h139 == _T_12323 ? _GEN_4 : mem_313;
  assign _GEN_8512 = 11'h13a == _T_12323 ? _GEN_4 : mem_314;
  assign _GEN_8513 = 11'h13b == _T_12323 ? _GEN_4 : mem_315;
  assign _GEN_8514 = 11'h13c == _T_12323 ? _GEN_4 : mem_316;
  assign _GEN_8515 = 11'h13d == _T_12323 ? _GEN_4 : mem_317;
  assign _GEN_8516 = 11'h13e == _T_12323 ? _GEN_4 : mem_318;
  assign _GEN_8517 = 11'h13f == _T_12323 ? _GEN_4 : mem_319;
  assign _GEN_8518 = 11'h140 == _T_12323 ? _GEN_4 : mem_320;
  assign _GEN_8519 = 11'h141 == _T_12323 ? _GEN_4 : mem_321;
  assign _GEN_8520 = 11'h142 == _T_12323 ? _GEN_4 : mem_322;
  assign _GEN_8521 = 11'h143 == _T_12323 ? _GEN_4 : mem_323;
  assign _GEN_8522 = 11'h144 == _T_12323 ? _GEN_4 : mem_324;
  assign _GEN_8523 = 11'h145 == _T_12323 ? _GEN_4 : mem_325;
  assign _GEN_8524 = 11'h146 == _T_12323 ? _GEN_4 : mem_326;
  assign _GEN_8525 = 11'h147 == _T_12323 ? _GEN_4 : mem_327;
  assign _GEN_8526 = 11'h148 == _T_12323 ? _GEN_4 : mem_328;
  assign _GEN_8527 = 11'h149 == _T_12323 ? _GEN_4 : mem_329;
  assign _GEN_8528 = 11'h14a == _T_12323 ? _GEN_4 : mem_330;
  assign _GEN_8529 = 11'h14b == _T_12323 ? _GEN_4 : mem_331;
  assign _GEN_8530 = 11'h14c == _T_12323 ? _GEN_4 : mem_332;
  assign _GEN_8531 = 11'h14d == _T_12323 ? _GEN_4 : mem_333;
  assign _GEN_8532 = 11'h14e == _T_12323 ? _GEN_4 : mem_334;
  assign _GEN_8533 = 11'h14f == _T_12323 ? _GEN_4 : mem_335;
  assign _GEN_8534 = 11'h150 == _T_12323 ? _GEN_4 : mem_336;
  assign _GEN_8535 = 11'h151 == _T_12323 ? _GEN_4 : mem_337;
  assign _GEN_8536 = 11'h152 == _T_12323 ? _GEN_4 : mem_338;
  assign _GEN_8537 = 11'h153 == _T_12323 ? _GEN_4 : mem_339;
  assign _GEN_8538 = 11'h154 == _T_12323 ? _GEN_4 : mem_340;
  assign _GEN_8539 = 11'h155 == _T_12323 ? _GEN_4 : mem_341;
  assign _GEN_8540 = 11'h156 == _T_12323 ? _GEN_4 : mem_342;
  assign _GEN_8541 = 11'h157 == _T_12323 ? _GEN_4 : mem_343;
  assign _GEN_8542 = 11'h158 == _T_12323 ? _GEN_4 : mem_344;
  assign _GEN_8543 = 11'h159 == _T_12323 ? _GEN_4 : mem_345;
  assign _GEN_8544 = 11'h15a == _T_12323 ? _GEN_4 : mem_346;
  assign _GEN_8545 = 11'h15b == _T_12323 ? _GEN_4 : mem_347;
  assign _GEN_8546 = 11'h15c == _T_12323 ? _GEN_4 : mem_348;
  assign _GEN_8547 = 11'h15d == _T_12323 ? _GEN_4 : mem_349;
  assign _GEN_8548 = 11'h15e == _T_12323 ? _GEN_4 : mem_350;
  assign _GEN_8549 = 11'h15f == _T_12323 ? _GEN_4 : mem_351;
  assign _GEN_8550 = 11'h160 == _T_12323 ? _GEN_4 : mem_352;
  assign _GEN_8551 = 11'h161 == _T_12323 ? _GEN_4 : mem_353;
  assign _GEN_8552 = 11'h162 == _T_12323 ? _GEN_4 : mem_354;
  assign _GEN_8553 = 11'h163 == _T_12323 ? _GEN_4 : mem_355;
  assign _GEN_8554 = 11'h164 == _T_12323 ? _GEN_4 : mem_356;
  assign _GEN_8555 = 11'h165 == _T_12323 ? _GEN_4 : mem_357;
  assign _GEN_8556 = 11'h166 == _T_12323 ? _GEN_4 : mem_358;
  assign _GEN_8557 = 11'h167 == _T_12323 ? _GEN_4 : mem_359;
  assign _GEN_8558 = 11'h168 == _T_12323 ? _GEN_4 : mem_360;
  assign _GEN_8559 = 11'h169 == _T_12323 ? _GEN_4 : mem_361;
  assign _GEN_8560 = 11'h16a == _T_12323 ? _GEN_4 : mem_362;
  assign _GEN_8561 = 11'h16b == _T_12323 ? _GEN_4 : mem_363;
  assign _GEN_8562 = 11'h16c == _T_12323 ? _GEN_4 : mem_364;
  assign _GEN_8563 = 11'h16d == _T_12323 ? _GEN_4 : mem_365;
  assign _GEN_8564 = 11'h16e == _T_12323 ? _GEN_4 : mem_366;
  assign _GEN_8565 = 11'h16f == _T_12323 ? _GEN_4 : mem_367;
  assign _GEN_8566 = 11'h170 == _T_12323 ? _GEN_4 : mem_368;
  assign _GEN_8567 = 11'h171 == _T_12323 ? _GEN_4 : mem_369;
  assign _GEN_8568 = 11'h172 == _T_12323 ? _GEN_4 : mem_370;
  assign _GEN_8569 = 11'h173 == _T_12323 ? _GEN_4 : mem_371;
  assign _GEN_8570 = 11'h174 == _T_12323 ? _GEN_4 : mem_372;
  assign _GEN_8571 = 11'h175 == _T_12323 ? _GEN_4 : mem_373;
  assign _GEN_8572 = 11'h176 == _T_12323 ? _GEN_4 : mem_374;
  assign _GEN_8573 = 11'h177 == _T_12323 ? _GEN_4 : mem_375;
  assign _GEN_8574 = 11'h178 == _T_12323 ? _GEN_4 : mem_376;
  assign _GEN_8575 = 11'h179 == _T_12323 ? _GEN_4 : mem_377;
  assign _GEN_8576 = 11'h17a == _T_12323 ? _GEN_4 : mem_378;
  assign _GEN_8577 = 11'h17b == _T_12323 ? _GEN_4 : mem_379;
  assign _GEN_8578 = 11'h17c == _T_12323 ? _GEN_4 : mem_380;
  assign _GEN_8579 = 11'h17d == _T_12323 ? _GEN_4 : mem_381;
  assign _GEN_8580 = 11'h17e == _T_12323 ? _GEN_4 : mem_382;
  assign _GEN_8581 = 11'h17f == _T_12323 ? _GEN_4 : mem_383;
  assign _GEN_8582 = 11'h180 == _T_12323 ? _GEN_4 : mem_384;
  assign _GEN_8583 = 11'h181 == _T_12323 ? _GEN_4 : mem_385;
  assign _GEN_8584 = 11'h182 == _T_12323 ? _GEN_4 : mem_386;
  assign _GEN_8585 = 11'h183 == _T_12323 ? _GEN_4 : mem_387;
  assign _GEN_8586 = 11'h184 == _T_12323 ? _GEN_4 : mem_388;
  assign _GEN_8587 = 11'h185 == _T_12323 ? _GEN_4 : mem_389;
  assign _GEN_8588 = 11'h186 == _T_12323 ? _GEN_4 : mem_390;
  assign _GEN_8589 = 11'h187 == _T_12323 ? _GEN_4 : mem_391;
  assign _GEN_8590 = 11'h188 == _T_12323 ? _GEN_4 : mem_392;
  assign _GEN_8591 = 11'h189 == _T_12323 ? _GEN_4 : mem_393;
  assign _GEN_8592 = 11'h18a == _T_12323 ? _GEN_4 : mem_394;
  assign _GEN_8593 = 11'h18b == _T_12323 ? _GEN_4 : mem_395;
  assign _GEN_8594 = 11'h18c == _T_12323 ? _GEN_4 : mem_396;
  assign _GEN_8595 = 11'h18d == _T_12323 ? _GEN_4 : mem_397;
  assign _GEN_8596 = 11'h18e == _T_12323 ? _GEN_4 : mem_398;
  assign _GEN_8597 = 11'h18f == _T_12323 ? _GEN_4 : mem_399;
  assign _GEN_8598 = 11'h190 == _T_12323 ? _GEN_4 : mem_400;
  assign _GEN_8599 = 11'h191 == _T_12323 ? _GEN_4 : mem_401;
  assign _GEN_8600 = 11'h192 == _T_12323 ? _GEN_4 : mem_402;
  assign _GEN_8601 = 11'h193 == _T_12323 ? _GEN_4 : mem_403;
  assign _GEN_8602 = 11'h194 == _T_12323 ? _GEN_4 : mem_404;
  assign _GEN_8603 = 11'h195 == _T_12323 ? _GEN_4 : mem_405;
  assign _GEN_8604 = 11'h196 == _T_12323 ? _GEN_4 : mem_406;
  assign _GEN_8605 = 11'h197 == _T_12323 ? _GEN_4 : mem_407;
  assign _GEN_8606 = 11'h198 == _T_12323 ? _GEN_4 : mem_408;
  assign _GEN_8607 = 11'h199 == _T_12323 ? _GEN_4 : mem_409;
  assign _GEN_8608 = 11'h19a == _T_12323 ? _GEN_4 : mem_410;
  assign _GEN_8609 = 11'h19b == _T_12323 ? _GEN_4 : mem_411;
  assign _GEN_8610 = 11'h19c == _T_12323 ? _GEN_4 : mem_412;
  assign _GEN_8611 = 11'h19d == _T_12323 ? _GEN_4 : mem_413;
  assign _GEN_8612 = 11'h19e == _T_12323 ? _GEN_4 : mem_414;
  assign _GEN_8613 = 11'h19f == _T_12323 ? _GEN_4 : mem_415;
  assign _GEN_8614 = 11'h1a0 == _T_12323 ? _GEN_4 : mem_416;
  assign _GEN_8615 = 11'h1a1 == _T_12323 ? _GEN_4 : mem_417;
  assign _GEN_8616 = 11'h1a2 == _T_12323 ? _GEN_4 : mem_418;
  assign _GEN_8617 = 11'h1a3 == _T_12323 ? _GEN_4 : mem_419;
  assign _GEN_8618 = 11'h1a4 == _T_12323 ? _GEN_4 : mem_420;
  assign _GEN_8619 = 11'h1a5 == _T_12323 ? _GEN_4 : mem_421;
  assign _GEN_8620 = 11'h1a6 == _T_12323 ? _GEN_4 : mem_422;
  assign _GEN_8621 = 11'h1a7 == _T_12323 ? _GEN_4 : mem_423;
  assign _GEN_8622 = 11'h1a8 == _T_12323 ? _GEN_4 : mem_424;
  assign _GEN_8623 = 11'h1a9 == _T_12323 ? _GEN_4 : mem_425;
  assign _GEN_8624 = 11'h1aa == _T_12323 ? _GEN_4 : mem_426;
  assign _GEN_8625 = 11'h1ab == _T_12323 ? _GEN_4 : mem_427;
  assign _GEN_8626 = 11'h1ac == _T_12323 ? _GEN_4 : mem_428;
  assign _GEN_8627 = 11'h1ad == _T_12323 ? _GEN_4 : mem_429;
  assign _GEN_8628 = 11'h1ae == _T_12323 ? _GEN_4 : mem_430;
  assign _GEN_8629 = 11'h1af == _T_12323 ? _GEN_4 : mem_431;
  assign _GEN_8630 = 11'h1b0 == _T_12323 ? _GEN_4 : mem_432;
  assign _GEN_8631 = 11'h1b1 == _T_12323 ? _GEN_4 : mem_433;
  assign _GEN_8632 = 11'h1b2 == _T_12323 ? _GEN_4 : mem_434;
  assign _GEN_8633 = 11'h1b3 == _T_12323 ? _GEN_4 : mem_435;
  assign _GEN_8634 = 11'h1b4 == _T_12323 ? _GEN_4 : mem_436;
  assign _GEN_8635 = 11'h1b5 == _T_12323 ? _GEN_4 : mem_437;
  assign _GEN_8636 = 11'h1b6 == _T_12323 ? _GEN_4 : mem_438;
  assign _GEN_8637 = 11'h1b7 == _T_12323 ? _GEN_4 : mem_439;
  assign _GEN_8638 = 11'h1b8 == _T_12323 ? _GEN_4 : mem_440;
  assign _GEN_8639 = 11'h1b9 == _T_12323 ? _GEN_4 : mem_441;
  assign _GEN_8640 = 11'h1ba == _T_12323 ? _GEN_4 : mem_442;
  assign _GEN_8641 = 11'h1bb == _T_12323 ? _GEN_4 : mem_443;
  assign _GEN_8642 = 11'h1bc == _T_12323 ? _GEN_4 : mem_444;
  assign _GEN_8643 = 11'h1bd == _T_12323 ? _GEN_4 : mem_445;
  assign _GEN_8644 = 11'h1be == _T_12323 ? _GEN_4 : mem_446;
  assign _GEN_8645 = 11'h1bf == _T_12323 ? _GEN_4 : mem_447;
  assign _GEN_8646 = 11'h1c0 == _T_12323 ? _GEN_4 : mem_448;
  assign _GEN_8647 = 11'h1c1 == _T_12323 ? _GEN_4 : mem_449;
  assign _GEN_8648 = 11'h1c2 == _T_12323 ? _GEN_4 : mem_450;
  assign _GEN_8649 = 11'h1c3 == _T_12323 ? _GEN_4 : mem_451;
  assign _GEN_8650 = 11'h1c4 == _T_12323 ? _GEN_4 : mem_452;
  assign _GEN_8651 = 11'h1c5 == _T_12323 ? _GEN_4 : mem_453;
  assign _GEN_8652 = 11'h1c6 == _T_12323 ? _GEN_4 : mem_454;
  assign _GEN_8653 = 11'h1c7 == _T_12323 ? _GEN_4 : mem_455;
  assign _GEN_8654 = 11'h1c8 == _T_12323 ? _GEN_4 : mem_456;
  assign _GEN_8655 = 11'h1c9 == _T_12323 ? _GEN_4 : mem_457;
  assign _GEN_8656 = 11'h1ca == _T_12323 ? _GEN_4 : mem_458;
  assign _GEN_8657 = 11'h1cb == _T_12323 ? _GEN_4 : mem_459;
  assign _GEN_8658 = 11'h1cc == _T_12323 ? _GEN_4 : mem_460;
  assign _GEN_8659 = 11'h1cd == _T_12323 ? _GEN_4 : mem_461;
  assign _GEN_8660 = 11'h1ce == _T_12323 ? _GEN_4 : mem_462;
  assign _GEN_8661 = 11'h1cf == _T_12323 ? _GEN_4 : mem_463;
  assign _GEN_8662 = 11'h1d0 == _T_12323 ? _GEN_4 : mem_464;
  assign _GEN_8663 = 11'h1d1 == _T_12323 ? _GEN_4 : mem_465;
  assign _GEN_8664 = 11'h1d2 == _T_12323 ? _GEN_4 : mem_466;
  assign _GEN_8665 = 11'h1d3 == _T_12323 ? _GEN_4 : mem_467;
  assign _GEN_8666 = 11'h1d4 == _T_12323 ? _GEN_4 : mem_468;
  assign _GEN_8667 = 11'h1d5 == _T_12323 ? _GEN_4 : mem_469;
  assign _GEN_8668 = 11'h1d6 == _T_12323 ? _GEN_4 : mem_470;
  assign _GEN_8669 = 11'h1d7 == _T_12323 ? _GEN_4 : mem_471;
  assign _GEN_8670 = 11'h1d8 == _T_12323 ? _GEN_4 : mem_472;
  assign _GEN_8671 = 11'h1d9 == _T_12323 ? _GEN_4 : mem_473;
  assign _GEN_8672 = 11'h1da == _T_12323 ? _GEN_4 : mem_474;
  assign _GEN_8673 = 11'h1db == _T_12323 ? _GEN_4 : mem_475;
  assign _GEN_8674 = 11'h1dc == _T_12323 ? _GEN_4 : mem_476;
  assign _GEN_8675 = 11'h1dd == _T_12323 ? _GEN_4 : mem_477;
  assign _GEN_8676 = 11'h1de == _T_12323 ? _GEN_4 : mem_478;
  assign _GEN_8677 = 11'h1df == _T_12323 ? _GEN_4 : mem_479;
  assign _GEN_8678 = 11'h1e0 == _T_12323 ? _GEN_4 : mem_480;
  assign _GEN_8679 = 11'h1e1 == _T_12323 ? _GEN_4 : mem_481;
  assign _GEN_8680 = 11'h1e2 == _T_12323 ? _GEN_4 : mem_482;
  assign _GEN_8681 = 11'h1e3 == _T_12323 ? _GEN_4 : mem_483;
  assign _GEN_8682 = 11'h1e4 == _T_12323 ? _GEN_4 : mem_484;
  assign _GEN_8683 = 11'h1e5 == _T_12323 ? _GEN_4 : mem_485;
  assign _GEN_8684 = 11'h1e6 == _T_12323 ? _GEN_4 : mem_486;
  assign _GEN_8685 = 11'h1e7 == _T_12323 ? _GEN_4 : mem_487;
  assign _GEN_8686 = 11'h1e8 == _T_12323 ? _GEN_4 : mem_488;
  assign _GEN_8687 = 11'h1e9 == _T_12323 ? _GEN_4 : mem_489;
  assign _GEN_8688 = 11'h1ea == _T_12323 ? _GEN_4 : mem_490;
  assign _GEN_8689 = 11'h1eb == _T_12323 ? _GEN_4 : mem_491;
  assign _GEN_8690 = 11'h1ec == _T_12323 ? _GEN_4 : mem_492;
  assign _GEN_8691 = 11'h1ed == _T_12323 ? _GEN_4 : mem_493;
  assign _GEN_8692 = 11'h1ee == _T_12323 ? _GEN_4 : mem_494;
  assign _GEN_8693 = 11'h1ef == _T_12323 ? _GEN_4 : mem_495;
  assign _GEN_8694 = 11'h1f0 == _T_12323 ? _GEN_4 : mem_496;
  assign _GEN_8695 = 11'h1f1 == _T_12323 ? _GEN_4 : mem_497;
  assign _GEN_8696 = 11'h1f2 == _T_12323 ? _GEN_4 : mem_498;
  assign _GEN_8697 = 11'h1f3 == _T_12323 ? _GEN_4 : mem_499;
  assign _GEN_8698 = 11'h1f4 == _T_12323 ? _GEN_4 : mem_500;
  assign _GEN_8699 = 11'h1f5 == _T_12323 ? _GEN_4 : mem_501;
  assign _GEN_8700 = 11'h1f6 == _T_12323 ? _GEN_4 : mem_502;
  assign _GEN_8701 = 11'h1f7 == _T_12323 ? _GEN_4 : mem_503;
  assign _GEN_8702 = 11'h1f8 == _T_12323 ? _GEN_4 : mem_504;
  assign _GEN_8703 = 11'h1f9 == _T_12323 ? _GEN_4 : mem_505;
  assign _GEN_8704 = 11'h1fa == _T_12323 ? _GEN_4 : mem_506;
  assign _GEN_8705 = 11'h1fb == _T_12323 ? _GEN_4 : mem_507;
  assign _GEN_8706 = 11'h1fc == _T_12323 ? _GEN_4 : mem_508;
  assign _GEN_8707 = 11'h1fd == _T_12323 ? _GEN_4 : mem_509;
  assign _GEN_8708 = 11'h1fe == _T_12323 ? _GEN_4 : mem_510;
  assign _GEN_8709 = 11'h1ff == _T_12323 ? _GEN_4 : mem_511;
  assign _GEN_8710 = 11'h200 == _T_12323 ? _GEN_4 : mem_512;
  assign _GEN_8711 = 11'h201 == _T_12323 ? _GEN_4 : mem_513;
  assign _GEN_8712 = 11'h202 == _T_12323 ? _GEN_4 : mem_514;
  assign _GEN_8713 = 11'h203 == _T_12323 ? _GEN_4 : mem_515;
  assign _GEN_8714 = 11'h204 == _T_12323 ? _GEN_4 : mem_516;
  assign _GEN_8715 = 11'h205 == _T_12323 ? _GEN_4 : mem_517;
  assign _GEN_8716 = 11'h206 == _T_12323 ? _GEN_4 : mem_518;
  assign _GEN_8717 = 11'h207 == _T_12323 ? _GEN_4 : mem_519;
  assign _GEN_8718 = 11'h208 == _T_12323 ? _GEN_4 : mem_520;
  assign _GEN_8719 = 11'h209 == _T_12323 ? _GEN_4 : mem_521;
  assign _GEN_8720 = 11'h20a == _T_12323 ? _GEN_4 : mem_522;
  assign _GEN_8721 = 11'h20b == _T_12323 ? _GEN_4 : mem_523;
  assign _GEN_8722 = 11'h20c == _T_12323 ? _GEN_4 : mem_524;
  assign _GEN_8723 = 11'h20d == _T_12323 ? _GEN_4 : mem_525;
  assign _GEN_8724 = 11'h20e == _T_12323 ? _GEN_4 : mem_526;
  assign _GEN_8725 = 11'h20f == _T_12323 ? _GEN_4 : mem_527;
  assign _GEN_8726 = 11'h210 == _T_12323 ? _GEN_4 : mem_528;
  assign _GEN_8727 = 11'h211 == _T_12323 ? _GEN_4 : mem_529;
  assign _GEN_8728 = 11'h212 == _T_12323 ? _GEN_4 : mem_530;
  assign _GEN_8729 = 11'h213 == _T_12323 ? _GEN_4 : mem_531;
  assign _GEN_8730 = 11'h214 == _T_12323 ? _GEN_4 : mem_532;
  assign _GEN_8731 = 11'h215 == _T_12323 ? _GEN_4 : mem_533;
  assign _GEN_8732 = 11'h216 == _T_12323 ? _GEN_4 : mem_534;
  assign _GEN_8733 = 11'h217 == _T_12323 ? _GEN_4 : mem_535;
  assign _GEN_8734 = 11'h218 == _T_12323 ? _GEN_4 : mem_536;
  assign _GEN_8735 = 11'h219 == _T_12323 ? _GEN_4 : mem_537;
  assign _GEN_8736 = 11'h21a == _T_12323 ? _GEN_4 : mem_538;
  assign _GEN_8737 = 11'h21b == _T_12323 ? _GEN_4 : mem_539;
  assign _GEN_8738 = 11'h21c == _T_12323 ? _GEN_4 : mem_540;
  assign _GEN_8739 = 11'h21d == _T_12323 ? _GEN_4 : mem_541;
  assign _GEN_8740 = 11'h21e == _T_12323 ? _GEN_4 : mem_542;
  assign _GEN_8741 = 11'h21f == _T_12323 ? _GEN_4 : mem_543;
  assign _GEN_8742 = 11'h220 == _T_12323 ? _GEN_4 : mem_544;
  assign _GEN_8743 = 11'h221 == _T_12323 ? _GEN_4 : mem_545;
  assign _GEN_8744 = 11'h222 == _T_12323 ? _GEN_4 : mem_546;
  assign _GEN_8745 = 11'h223 == _T_12323 ? _GEN_4 : mem_547;
  assign _GEN_8746 = 11'h224 == _T_12323 ? _GEN_4 : mem_548;
  assign _GEN_8747 = 11'h225 == _T_12323 ? _GEN_4 : mem_549;
  assign _GEN_8748 = 11'h226 == _T_12323 ? _GEN_4 : mem_550;
  assign _GEN_8749 = 11'h227 == _T_12323 ? _GEN_4 : mem_551;
  assign _GEN_8750 = 11'h228 == _T_12323 ? _GEN_4 : mem_552;
  assign _GEN_8751 = 11'h229 == _T_12323 ? _GEN_4 : mem_553;
  assign _GEN_8752 = 11'h22a == _T_12323 ? _GEN_4 : mem_554;
  assign _GEN_8753 = 11'h22b == _T_12323 ? _GEN_4 : mem_555;
  assign _GEN_8754 = 11'h22c == _T_12323 ? _GEN_4 : mem_556;
  assign _GEN_8755 = 11'h22d == _T_12323 ? _GEN_4 : mem_557;
  assign _GEN_8756 = 11'h22e == _T_12323 ? _GEN_4 : mem_558;
  assign _GEN_8757 = 11'h22f == _T_12323 ? _GEN_4 : mem_559;
  assign _GEN_8758 = 11'h230 == _T_12323 ? _GEN_4 : mem_560;
  assign _GEN_8759 = 11'h231 == _T_12323 ? _GEN_4 : mem_561;
  assign _GEN_8760 = 11'h232 == _T_12323 ? _GEN_4 : mem_562;
  assign _GEN_8761 = 11'h233 == _T_12323 ? _GEN_4 : mem_563;
  assign _GEN_8762 = 11'h234 == _T_12323 ? _GEN_4 : mem_564;
  assign _GEN_8763 = 11'h235 == _T_12323 ? _GEN_4 : mem_565;
  assign _GEN_8764 = 11'h236 == _T_12323 ? _GEN_4 : mem_566;
  assign _GEN_8765 = 11'h237 == _T_12323 ? _GEN_4 : mem_567;
  assign _GEN_8766 = 11'h238 == _T_12323 ? _GEN_4 : mem_568;
  assign _GEN_8767 = 11'h239 == _T_12323 ? _GEN_4 : mem_569;
  assign _GEN_8768 = 11'h23a == _T_12323 ? _GEN_4 : mem_570;
  assign _GEN_8769 = 11'h23b == _T_12323 ? _GEN_4 : mem_571;
  assign _GEN_8770 = 11'h23c == _T_12323 ? _GEN_4 : mem_572;
  assign _GEN_8771 = 11'h23d == _T_12323 ? _GEN_4 : mem_573;
  assign _GEN_8772 = 11'h23e == _T_12323 ? _GEN_4 : mem_574;
  assign _GEN_8773 = 11'h23f == _T_12323 ? _GEN_4 : mem_575;
  assign _GEN_8774 = 11'h240 == _T_12323 ? _GEN_4 : mem_576;
  assign _GEN_8775 = 11'h241 == _T_12323 ? _GEN_4 : mem_577;
  assign _GEN_8776 = 11'h242 == _T_12323 ? _GEN_4 : mem_578;
  assign _GEN_8777 = 11'h243 == _T_12323 ? _GEN_4 : mem_579;
  assign _GEN_8778 = 11'h244 == _T_12323 ? _GEN_4 : mem_580;
  assign _GEN_8779 = 11'h245 == _T_12323 ? _GEN_4 : mem_581;
  assign _GEN_8780 = 11'h246 == _T_12323 ? _GEN_4 : mem_582;
  assign _GEN_8781 = 11'h247 == _T_12323 ? _GEN_4 : mem_583;
  assign _GEN_8782 = 11'h248 == _T_12323 ? _GEN_4 : mem_584;
  assign _GEN_8783 = 11'h249 == _T_12323 ? _GEN_4 : mem_585;
  assign _GEN_8784 = 11'h24a == _T_12323 ? _GEN_4 : mem_586;
  assign _GEN_8785 = 11'h24b == _T_12323 ? _GEN_4 : mem_587;
  assign _GEN_8786 = 11'h24c == _T_12323 ? _GEN_4 : mem_588;
  assign _GEN_8787 = 11'h24d == _T_12323 ? _GEN_4 : mem_589;
  assign _GEN_8788 = 11'h24e == _T_12323 ? _GEN_4 : mem_590;
  assign _GEN_8789 = 11'h24f == _T_12323 ? _GEN_4 : mem_591;
  assign _GEN_8790 = 11'h250 == _T_12323 ? _GEN_4 : mem_592;
  assign _GEN_8791 = 11'h251 == _T_12323 ? _GEN_4 : mem_593;
  assign _GEN_8792 = 11'h252 == _T_12323 ? _GEN_4 : mem_594;
  assign _GEN_8793 = 11'h253 == _T_12323 ? _GEN_4 : mem_595;
  assign _GEN_8794 = 11'h254 == _T_12323 ? _GEN_4 : mem_596;
  assign _GEN_8795 = 11'h255 == _T_12323 ? _GEN_4 : mem_597;
  assign _GEN_8796 = 11'h256 == _T_12323 ? _GEN_4 : mem_598;
  assign _GEN_8797 = 11'h257 == _T_12323 ? _GEN_4 : mem_599;
  assign _GEN_8798 = 11'h258 == _T_12323 ? _GEN_4 : mem_600;
  assign _GEN_8799 = 11'h259 == _T_12323 ? _GEN_4 : mem_601;
  assign _GEN_8800 = 11'h25a == _T_12323 ? _GEN_4 : mem_602;
  assign _GEN_8801 = 11'h25b == _T_12323 ? _GEN_4 : mem_603;
  assign _GEN_8802 = 11'h25c == _T_12323 ? _GEN_4 : mem_604;
  assign _GEN_8803 = 11'h25d == _T_12323 ? _GEN_4 : mem_605;
  assign _GEN_8804 = 11'h25e == _T_12323 ? _GEN_4 : mem_606;
  assign _GEN_8805 = 11'h25f == _T_12323 ? _GEN_4 : mem_607;
  assign _GEN_8806 = 11'h260 == _T_12323 ? _GEN_4 : mem_608;
  assign _GEN_8807 = 11'h261 == _T_12323 ? _GEN_4 : mem_609;
  assign _GEN_8808 = 11'h262 == _T_12323 ? _GEN_4 : mem_610;
  assign _GEN_8809 = 11'h263 == _T_12323 ? _GEN_4 : mem_611;
  assign _GEN_8810 = 11'h264 == _T_12323 ? _GEN_4 : mem_612;
  assign _GEN_8811 = 11'h265 == _T_12323 ? _GEN_4 : mem_613;
  assign _GEN_8812 = 11'h266 == _T_12323 ? _GEN_4 : mem_614;
  assign _GEN_8813 = 11'h267 == _T_12323 ? _GEN_4 : mem_615;
  assign _GEN_8814 = 11'h268 == _T_12323 ? _GEN_4 : mem_616;
  assign _GEN_8815 = 11'h269 == _T_12323 ? _GEN_4 : mem_617;
  assign _GEN_8816 = 11'h26a == _T_12323 ? _GEN_4 : mem_618;
  assign _GEN_8817 = 11'h26b == _T_12323 ? _GEN_4 : mem_619;
  assign _GEN_8818 = 11'h26c == _T_12323 ? _GEN_4 : mem_620;
  assign _GEN_8819 = 11'h26d == _T_12323 ? _GEN_4 : mem_621;
  assign _GEN_8820 = 11'h26e == _T_12323 ? _GEN_4 : mem_622;
  assign _GEN_8821 = 11'h26f == _T_12323 ? _GEN_4 : mem_623;
  assign _GEN_8822 = 11'h270 == _T_12323 ? _GEN_4 : mem_624;
  assign _GEN_8823 = 11'h271 == _T_12323 ? _GEN_4 : mem_625;
  assign _GEN_8824 = 11'h272 == _T_12323 ? _GEN_4 : mem_626;
  assign _GEN_8825 = 11'h273 == _T_12323 ? _GEN_4 : mem_627;
  assign _GEN_8826 = 11'h274 == _T_12323 ? _GEN_4 : mem_628;
  assign _GEN_8827 = 11'h275 == _T_12323 ? _GEN_4 : mem_629;
  assign _GEN_8828 = 11'h276 == _T_12323 ? _GEN_4 : mem_630;
  assign _GEN_8829 = 11'h277 == _T_12323 ? _GEN_4 : mem_631;
  assign _GEN_8830 = 11'h278 == _T_12323 ? _GEN_4 : mem_632;
  assign _GEN_8831 = 11'h279 == _T_12323 ? _GEN_4 : mem_633;
  assign _GEN_8832 = 11'h27a == _T_12323 ? _GEN_4 : mem_634;
  assign _GEN_8833 = 11'h27b == _T_12323 ? _GEN_4 : mem_635;
  assign _GEN_8834 = 11'h27c == _T_12323 ? _GEN_4 : mem_636;
  assign _GEN_8835 = 11'h27d == _T_12323 ? _GEN_4 : mem_637;
  assign _GEN_8836 = 11'h27e == _T_12323 ? _GEN_4 : mem_638;
  assign _GEN_8837 = 11'h27f == _T_12323 ? _GEN_4 : mem_639;
  assign _GEN_8838 = 11'h280 == _T_12323 ? _GEN_4 : mem_640;
  assign _GEN_8839 = 11'h281 == _T_12323 ? _GEN_4 : mem_641;
  assign _GEN_8840 = 11'h282 == _T_12323 ? _GEN_4 : mem_642;
  assign _GEN_8841 = 11'h283 == _T_12323 ? _GEN_4 : mem_643;
  assign _GEN_8842 = 11'h284 == _T_12323 ? _GEN_4 : mem_644;
  assign _GEN_8843 = 11'h285 == _T_12323 ? _GEN_4 : mem_645;
  assign _GEN_8844 = 11'h286 == _T_12323 ? _GEN_4 : mem_646;
  assign _GEN_8845 = 11'h287 == _T_12323 ? _GEN_4 : mem_647;
  assign _GEN_8846 = 11'h288 == _T_12323 ? _GEN_4 : mem_648;
  assign _GEN_8847 = 11'h289 == _T_12323 ? _GEN_4 : mem_649;
  assign _GEN_8848 = 11'h28a == _T_12323 ? _GEN_4 : mem_650;
  assign _GEN_8849 = 11'h28b == _T_12323 ? _GEN_4 : mem_651;
  assign _GEN_8850 = 11'h28c == _T_12323 ? _GEN_4 : mem_652;
  assign _GEN_8851 = 11'h28d == _T_12323 ? _GEN_4 : mem_653;
  assign _GEN_8852 = 11'h28e == _T_12323 ? _GEN_4 : mem_654;
  assign _GEN_8853 = 11'h28f == _T_12323 ? _GEN_4 : mem_655;
  assign _GEN_8854 = 11'h290 == _T_12323 ? _GEN_4 : mem_656;
  assign _GEN_8855 = 11'h291 == _T_12323 ? _GEN_4 : mem_657;
  assign _GEN_8856 = 11'h292 == _T_12323 ? _GEN_4 : mem_658;
  assign _GEN_8857 = 11'h293 == _T_12323 ? _GEN_4 : mem_659;
  assign _GEN_8858 = 11'h294 == _T_12323 ? _GEN_4 : mem_660;
  assign _GEN_8859 = 11'h295 == _T_12323 ? _GEN_4 : mem_661;
  assign _GEN_8860 = 11'h296 == _T_12323 ? _GEN_4 : mem_662;
  assign _GEN_8861 = 11'h297 == _T_12323 ? _GEN_4 : mem_663;
  assign _GEN_8862 = 11'h298 == _T_12323 ? _GEN_4 : mem_664;
  assign _GEN_8863 = 11'h299 == _T_12323 ? _GEN_4 : mem_665;
  assign _GEN_8864 = 11'h29a == _T_12323 ? _GEN_4 : mem_666;
  assign _GEN_8865 = 11'h29b == _T_12323 ? _GEN_4 : mem_667;
  assign _GEN_8866 = 11'h29c == _T_12323 ? _GEN_4 : mem_668;
  assign _GEN_8867 = 11'h29d == _T_12323 ? _GEN_4 : mem_669;
  assign _GEN_8868 = 11'h29e == _T_12323 ? _GEN_4 : mem_670;
  assign _GEN_8869 = 11'h29f == _T_12323 ? _GEN_4 : mem_671;
  assign _GEN_8870 = 11'h2a0 == _T_12323 ? _GEN_4 : mem_672;
  assign _GEN_8871 = 11'h2a1 == _T_12323 ? _GEN_4 : mem_673;
  assign _GEN_8872 = 11'h2a2 == _T_12323 ? _GEN_4 : mem_674;
  assign _GEN_8873 = 11'h2a3 == _T_12323 ? _GEN_4 : mem_675;
  assign _GEN_8874 = 11'h2a4 == _T_12323 ? _GEN_4 : mem_676;
  assign _GEN_8875 = 11'h2a5 == _T_12323 ? _GEN_4 : mem_677;
  assign _GEN_8876 = 11'h2a6 == _T_12323 ? _GEN_4 : mem_678;
  assign _GEN_8877 = 11'h2a7 == _T_12323 ? _GEN_4 : mem_679;
  assign _GEN_8878 = 11'h2a8 == _T_12323 ? _GEN_4 : mem_680;
  assign _GEN_8879 = 11'h2a9 == _T_12323 ? _GEN_4 : mem_681;
  assign _GEN_8880 = 11'h2aa == _T_12323 ? _GEN_4 : mem_682;
  assign _GEN_8881 = 11'h2ab == _T_12323 ? _GEN_4 : mem_683;
  assign _GEN_8882 = 11'h2ac == _T_12323 ? _GEN_4 : mem_684;
  assign _GEN_8883 = 11'h2ad == _T_12323 ? _GEN_4 : mem_685;
  assign _GEN_8884 = 11'h2ae == _T_12323 ? _GEN_4 : mem_686;
  assign _GEN_8885 = 11'h2af == _T_12323 ? _GEN_4 : mem_687;
  assign _GEN_8886 = 11'h2b0 == _T_12323 ? _GEN_4 : mem_688;
  assign _GEN_8887 = 11'h2b1 == _T_12323 ? _GEN_4 : mem_689;
  assign _GEN_8888 = 11'h2b2 == _T_12323 ? _GEN_4 : mem_690;
  assign _GEN_8889 = 11'h2b3 == _T_12323 ? _GEN_4 : mem_691;
  assign _GEN_8890 = 11'h2b4 == _T_12323 ? _GEN_4 : mem_692;
  assign _GEN_8891 = 11'h2b5 == _T_12323 ? _GEN_4 : mem_693;
  assign _GEN_8892 = 11'h2b6 == _T_12323 ? _GEN_4 : mem_694;
  assign _GEN_8893 = 11'h2b7 == _T_12323 ? _GEN_4 : mem_695;
  assign _GEN_8894 = 11'h2b8 == _T_12323 ? _GEN_4 : mem_696;
  assign _GEN_8895 = 11'h2b9 == _T_12323 ? _GEN_4 : mem_697;
  assign _GEN_8896 = 11'h2ba == _T_12323 ? _GEN_4 : mem_698;
  assign _GEN_8897 = 11'h2bb == _T_12323 ? _GEN_4 : mem_699;
  assign _GEN_8898 = 11'h2bc == _T_12323 ? _GEN_4 : mem_700;
  assign _GEN_8899 = 11'h2bd == _T_12323 ? _GEN_4 : mem_701;
  assign _GEN_8900 = 11'h2be == _T_12323 ? _GEN_4 : mem_702;
  assign _GEN_8901 = 11'h2bf == _T_12323 ? _GEN_4 : mem_703;
  assign _GEN_8902 = 11'h2c0 == _T_12323 ? _GEN_4 : mem_704;
  assign _GEN_8903 = 11'h2c1 == _T_12323 ? _GEN_4 : mem_705;
  assign _GEN_8904 = 11'h2c2 == _T_12323 ? _GEN_4 : mem_706;
  assign _GEN_8905 = 11'h2c3 == _T_12323 ? _GEN_4 : mem_707;
  assign _GEN_8906 = 11'h2c4 == _T_12323 ? _GEN_4 : mem_708;
  assign _GEN_8907 = 11'h2c5 == _T_12323 ? _GEN_4 : mem_709;
  assign _GEN_8908 = 11'h2c6 == _T_12323 ? _GEN_4 : mem_710;
  assign _GEN_8909 = 11'h2c7 == _T_12323 ? _GEN_4 : mem_711;
  assign _GEN_8910 = 11'h2c8 == _T_12323 ? _GEN_4 : mem_712;
  assign _GEN_8911 = 11'h2c9 == _T_12323 ? _GEN_4 : mem_713;
  assign _GEN_8912 = 11'h2ca == _T_12323 ? _GEN_4 : mem_714;
  assign _GEN_8913 = 11'h2cb == _T_12323 ? _GEN_4 : mem_715;
  assign _GEN_8914 = 11'h2cc == _T_12323 ? _GEN_4 : mem_716;
  assign _GEN_8915 = 11'h2cd == _T_12323 ? _GEN_4 : mem_717;
  assign _GEN_8916 = 11'h2ce == _T_12323 ? _GEN_4 : mem_718;
  assign _GEN_8917 = 11'h2cf == _T_12323 ? _GEN_4 : mem_719;
  assign _GEN_8918 = 11'h2d0 == _T_12323 ? _GEN_4 : mem_720;
  assign _GEN_8919 = 11'h2d1 == _T_12323 ? _GEN_4 : mem_721;
  assign _GEN_8920 = 11'h2d2 == _T_12323 ? _GEN_4 : mem_722;
  assign _GEN_8921 = 11'h2d3 == _T_12323 ? _GEN_4 : mem_723;
  assign _GEN_8922 = 11'h2d4 == _T_12323 ? _GEN_4 : mem_724;
  assign _GEN_8923 = 11'h2d5 == _T_12323 ? _GEN_4 : mem_725;
  assign _GEN_8924 = 11'h2d6 == _T_12323 ? _GEN_4 : mem_726;
  assign _GEN_8925 = 11'h2d7 == _T_12323 ? _GEN_4 : mem_727;
  assign _GEN_8926 = 11'h2d8 == _T_12323 ? _GEN_4 : mem_728;
  assign _GEN_8927 = 11'h2d9 == _T_12323 ? _GEN_4 : mem_729;
  assign _GEN_8928 = 11'h2da == _T_12323 ? _GEN_4 : mem_730;
  assign _GEN_8929 = 11'h2db == _T_12323 ? _GEN_4 : mem_731;
  assign _GEN_8930 = 11'h2dc == _T_12323 ? _GEN_4 : mem_732;
  assign _GEN_8931 = 11'h2dd == _T_12323 ? _GEN_4 : mem_733;
  assign _GEN_8932 = 11'h2de == _T_12323 ? _GEN_4 : mem_734;
  assign _GEN_8933 = 11'h2df == _T_12323 ? _GEN_4 : mem_735;
  assign _GEN_8934 = 11'h2e0 == _T_12323 ? _GEN_4 : mem_736;
  assign _GEN_8935 = 11'h2e1 == _T_12323 ? _GEN_4 : mem_737;
  assign _GEN_8936 = 11'h2e2 == _T_12323 ? _GEN_4 : mem_738;
  assign _GEN_8937 = 11'h2e3 == _T_12323 ? _GEN_4 : mem_739;
  assign _GEN_8938 = 11'h2e4 == _T_12323 ? _GEN_4 : mem_740;
  assign _GEN_8939 = 11'h2e5 == _T_12323 ? _GEN_4 : mem_741;
  assign _GEN_8940 = 11'h2e6 == _T_12323 ? _GEN_4 : mem_742;
  assign _GEN_8941 = 11'h2e7 == _T_12323 ? _GEN_4 : mem_743;
  assign _GEN_8942 = 11'h2e8 == _T_12323 ? _GEN_4 : mem_744;
  assign _GEN_8943 = 11'h2e9 == _T_12323 ? _GEN_4 : mem_745;
  assign _GEN_8944 = 11'h2ea == _T_12323 ? _GEN_4 : mem_746;
  assign _GEN_8945 = 11'h2eb == _T_12323 ? _GEN_4 : mem_747;
  assign _GEN_8946 = 11'h2ec == _T_12323 ? _GEN_4 : mem_748;
  assign _GEN_8947 = 11'h2ed == _T_12323 ? _GEN_4 : mem_749;
  assign _GEN_8948 = 11'h2ee == _T_12323 ? _GEN_4 : mem_750;
  assign _GEN_8949 = 11'h2ef == _T_12323 ? _GEN_4 : mem_751;
  assign _GEN_8950 = 11'h2f0 == _T_12323 ? _GEN_4 : mem_752;
  assign _GEN_8951 = 11'h2f1 == _T_12323 ? _GEN_4 : mem_753;
  assign _GEN_8952 = 11'h2f2 == _T_12323 ? _GEN_4 : mem_754;
  assign _GEN_8953 = 11'h2f3 == _T_12323 ? _GEN_4 : mem_755;
  assign _GEN_8954 = 11'h2f4 == _T_12323 ? _GEN_4 : mem_756;
  assign _GEN_8955 = 11'h2f5 == _T_12323 ? _GEN_4 : mem_757;
  assign _GEN_8956 = 11'h2f6 == _T_12323 ? _GEN_4 : mem_758;
  assign _GEN_8957 = 11'h2f7 == _T_12323 ? _GEN_4 : mem_759;
  assign _GEN_8958 = 11'h2f8 == _T_12323 ? _GEN_4 : mem_760;
  assign _GEN_8959 = 11'h2f9 == _T_12323 ? _GEN_4 : mem_761;
  assign _GEN_8960 = 11'h2fa == _T_12323 ? _GEN_4 : mem_762;
  assign _GEN_8961 = 11'h2fb == _T_12323 ? _GEN_4 : mem_763;
  assign _GEN_8962 = 11'h2fc == _T_12323 ? _GEN_4 : mem_764;
  assign _GEN_8963 = 11'h2fd == _T_12323 ? _GEN_4 : mem_765;
  assign _GEN_8964 = 11'h2fe == _T_12323 ? _GEN_4 : mem_766;
  assign _GEN_8965 = 11'h2ff == _T_12323 ? _GEN_4 : mem_767;
  assign _GEN_8966 = 11'h300 == _T_12323 ? _GEN_4 : mem_768;
  assign _GEN_8967 = 11'h301 == _T_12323 ? _GEN_4 : mem_769;
  assign _GEN_8968 = 11'h302 == _T_12323 ? _GEN_4 : mem_770;
  assign _GEN_8969 = 11'h303 == _T_12323 ? _GEN_4 : mem_771;
  assign _GEN_8970 = 11'h304 == _T_12323 ? _GEN_4 : mem_772;
  assign _GEN_8971 = 11'h305 == _T_12323 ? _GEN_4 : mem_773;
  assign _GEN_8972 = 11'h306 == _T_12323 ? _GEN_4 : mem_774;
  assign _GEN_8973 = 11'h307 == _T_12323 ? _GEN_4 : mem_775;
  assign _GEN_8974 = 11'h308 == _T_12323 ? _GEN_4 : mem_776;
  assign _GEN_8975 = 11'h309 == _T_12323 ? _GEN_4 : mem_777;
  assign _GEN_8976 = 11'h30a == _T_12323 ? _GEN_4 : mem_778;
  assign _GEN_8977 = 11'h30b == _T_12323 ? _GEN_4 : mem_779;
  assign _GEN_8978 = 11'h30c == _T_12323 ? _GEN_4 : mem_780;
  assign _GEN_8979 = 11'h30d == _T_12323 ? _GEN_4 : mem_781;
  assign _GEN_8980 = 11'h30e == _T_12323 ? _GEN_4 : mem_782;
  assign _GEN_8981 = 11'h30f == _T_12323 ? _GEN_4 : mem_783;
  assign _GEN_8982 = 11'h310 == _T_12323 ? _GEN_4 : mem_784;
  assign _GEN_8983 = 11'h311 == _T_12323 ? _GEN_4 : mem_785;
  assign _GEN_8984 = 11'h312 == _T_12323 ? _GEN_4 : mem_786;
  assign _GEN_8985 = 11'h313 == _T_12323 ? _GEN_4 : mem_787;
  assign _GEN_8986 = 11'h314 == _T_12323 ? _GEN_4 : mem_788;
  assign _GEN_8987 = 11'h315 == _T_12323 ? _GEN_4 : mem_789;
  assign _GEN_8988 = 11'h316 == _T_12323 ? _GEN_4 : mem_790;
  assign _GEN_8989 = 11'h317 == _T_12323 ? _GEN_4 : mem_791;
  assign _GEN_8990 = 11'h318 == _T_12323 ? _GEN_4 : mem_792;
  assign _GEN_8991 = 11'h319 == _T_12323 ? _GEN_4 : mem_793;
  assign _GEN_8992 = 11'h31a == _T_12323 ? _GEN_4 : mem_794;
  assign _GEN_8993 = 11'h31b == _T_12323 ? _GEN_4 : mem_795;
  assign _GEN_8994 = 11'h31c == _T_12323 ? _GEN_4 : mem_796;
  assign _GEN_8995 = 11'h31d == _T_12323 ? _GEN_4 : mem_797;
  assign _GEN_8996 = 11'h31e == _T_12323 ? _GEN_4 : mem_798;
  assign _GEN_8997 = 11'h31f == _T_12323 ? _GEN_4 : mem_799;
  assign _GEN_8998 = 11'h320 == _T_12323 ? _GEN_4 : mem_800;
  assign _GEN_8999 = 11'h321 == _T_12323 ? _GEN_4 : mem_801;
  assign _GEN_9000 = 11'h322 == _T_12323 ? _GEN_4 : mem_802;
  assign _GEN_9001 = 11'h323 == _T_12323 ? _GEN_4 : mem_803;
  assign _GEN_9002 = 11'h324 == _T_12323 ? _GEN_4 : mem_804;
  assign _GEN_9003 = 11'h325 == _T_12323 ? _GEN_4 : mem_805;
  assign _GEN_9004 = 11'h326 == _T_12323 ? _GEN_4 : mem_806;
  assign _GEN_9005 = 11'h327 == _T_12323 ? _GEN_4 : mem_807;
  assign _GEN_9006 = 11'h328 == _T_12323 ? _GEN_4 : mem_808;
  assign _GEN_9007 = 11'h329 == _T_12323 ? _GEN_4 : mem_809;
  assign _GEN_9008 = 11'h32a == _T_12323 ? _GEN_4 : mem_810;
  assign _GEN_9009 = 11'h32b == _T_12323 ? _GEN_4 : mem_811;
  assign _GEN_9010 = 11'h32c == _T_12323 ? _GEN_4 : mem_812;
  assign _GEN_9011 = 11'h32d == _T_12323 ? _GEN_4 : mem_813;
  assign _GEN_9012 = 11'h32e == _T_12323 ? _GEN_4 : mem_814;
  assign _GEN_9013 = 11'h32f == _T_12323 ? _GEN_4 : mem_815;
  assign _GEN_9014 = 11'h330 == _T_12323 ? _GEN_4 : mem_816;
  assign _GEN_9015 = 11'h331 == _T_12323 ? _GEN_4 : mem_817;
  assign _GEN_9016 = 11'h332 == _T_12323 ? _GEN_4 : mem_818;
  assign _GEN_9017 = 11'h333 == _T_12323 ? _GEN_4 : mem_819;
  assign _GEN_9018 = 11'h334 == _T_12323 ? _GEN_4 : mem_820;
  assign _GEN_9019 = 11'h335 == _T_12323 ? _GEN_4 : mem_821;
  assign _GEN_9020 = 11'h336 == _T_12323 ? _GEN_4 : mem_822;
  assign _GEN_9021 = 11'h337 == _T_12323 ? _GEN_4 : mem_823;
  assign _GEN_9022 = 11'h338 == _T_12323 ? _GEN_4 : mem_824;
  assign _GEN_9023 = 11'h339 == _T_12323 ? _GEN_4 : mem_825;
  assign _GEN_9024 = 11'h33a == _T_12323 ? _GEN_4 : mem_826;
  assign _GEN_9025 = 11'h33b == _T_12323 ? _GEN_4 : mem_827;
  assign _GEN_9026 = 11'h33c == _T_12323 ? _GEN_4 : mem_828;
  assign _GEN_9027 = 11'h33d == _T_12323 ? _GEN_4 : mem_829;
  assign _GEN_9028 = 11'h33e == _T_12323 ? _GEN_4 : mem_830;
  assign _GEN_9029 = 11'h33f == _T_12323 ? _GEN_4 : mem_831;
  assign _GEN_9030 = 11'h340 == _T_12323 ? _GEN_4 : mem_832;
  assign _GEN_9031 = 11'h341 == _T_12323 ? _GEN_4 : mem_833;
  assign _GEN_9032 = 11'h342 == _T_12323 ? _GEN_4 : mem_834;
  assign _GEN_9033 = 11'h343 == _T_12323 ? _GEN_4 : mem_835;
  assign _GEN_9034 = 11'h344 == _T_12323 ? _GEN_4 : mem_836;
  assign _GEN_9035 = 11'h345 == _T_12323 ? _GEN_4 : mem_837;
  assign _GEN_9036 = 11'h346 == _T_12323 ? _GEN_4 : mem_838;
  assign _GEN_9037 = 11'h347 == _T_12323 ? _GEN_4 : mem_839;
  assign _GEN_9038 = 11'h348 == _T_12323 ? _GEN_4 : mem_840;
  assign _GEN_9039 = 11'h349 == _T_12323 ? _GEN_4 : mem_841;
  assign _GEN_9040 = 11'h34a == _T_12323 ? _GEN_4 : mem_842;
  assign _GEN_9041 = 11'h34b == _T_12323 ? _GEN_4 : mem_843;
  assign _GEN_9042 = 11'h34c == _T_12323 ? _GEN_4 : mem_844;
  assign _GEN_9043 = 11'h34d == _T_12323 ? _GEN_4 : mem_845;
  assign _GEN_9044 = 11'h34e == _T_12323 ? _GEN_4 : mem_846;
  assign _GEN_9045 = 11'h34f == _T_12323 ? _GEN_4 : mem_847;
  assign _GEN_9046 = 11'h350 == _T_12323 ? _GEN_4 : mem_848;
  assign _GEN_9047 = 11'h351 == _T_12323 ? _GEN_4 : mem_849;
  assign _GEN_9048 = 11'h352 == _T_12323 ? _GEN_4 : mem_850;
  assign _GEN_9049 = 11'h353 == _T_12323 ? _GEN_4 : mem_851;
  assign _GEN_9050 = 11'h354 == _T_12323 ? _GEN_4 : mem_852;
  assign _GEN_9051 = 11'h355 == _T_12323 ? _GEN_4 : mem_853;
  assign _GEN_9052 = 11'h356 == _T_12323 ? _GEN_4 : mem_854;
  assign _GEN_9053 = 11'h357 == _T_12323 ? _GEN_4 : mem_855;
  assign _GEN_9054 = 11'h358 == _T_12323 ? _GEN_4 : mem_856;
  assign _GEN_9055 = 11'h359 == _T_12323 ? _GEN_4 : mem_857;
  assign _GEN_9056 = 11'h35a == _T_12323 ? _GEN_4 : mem_858;
  assign _GEN_9057 = 11'h35b == _T_12323 ? _GEN_4 : mem_859;
  assign _GEN_9058 = 11'h35c == _T_12323 ? _GEN_4 : mem_860;
  assign _GEN_9059 = 11'h35d == _T_12323 ? _GEN_4 : mem_861;
  assign _GEN_9060 = 11'h35e == _T_12323 ? _GEN_4 : mem_862;
  assign _GEN_9061 = 11'h35f == _T_12323 ? _GEN_4 : mem_863;
  assign _GEN_9062 = 11'h360 == _T_12323 ? _GEN_4 : mem_864;
  assign _GEN_9063 = 11'h361 == _T_12323 ? _GEN_4 : mem_865;
  assign _GEN_9064 = 11'h362 == _T_12323 ? _GEN_4 : mem_866;
  assign _GEN_9065 = 11'h363 == _T_12323 ? _GEN_4 : mem_867;
  assign _GEN_9066 = 11'h364 == _T_12323 ? _GEN_4 : mem_868;
  assign _GEN_9067 = 11'h365 == _T_12323 ? _GEN_4 : mem_869;
  assign _GEN_9068 = 11'h366 == _T_12323 ? _GEN_4 : mem_870;
  assign _GEN_9069 = 11'h367 == _T_12323 ? _GEN_4 : mem_871;
  assign _GEN_9070 = 11'h368 == _T_12323 ? _GEN_4 : mem_872;
  assign _GEN_9071 = 11'h369 == _T_12323 ? _GEN_4 : mem_873;
  assign _GEN_9072 = 11'h36a == _T_12323 ? _GEN_4 : mem_874;
  assign _GEN_9073 = 11'h36b == _T_12323 ? _GEN_4 : mem_875;
  assign _GEN_9074 = 11'h36c == _T_12323 ? _GEN_4 : mem_876;
  assign _GEN_9075 = 11'h36d == _T_12323 ? _GEN_4 : mem_877;
  assign _GEN_9076 = 11'h36e == _T_12323 ? _GEN_4 : mem_878;
  assign _GEN_9077 = 11'h36f == _T_12323 ? _GEN_4 : mem_879;
  assign _GEN_9078 = 11'h370 == _T_12323 ? _GEN_4 : mem_880;
  assign _GEN_9079 = 11'h371 == _T_12323 ? _GEN_4 : mem_881;
  assign _GEN_9080 = 11'h372 == _T_12323 ? _GEN_4 : mem_882;
  assign _GEN_9081 = 11'h373 == _T_12323 ? _GEN_4 : mem_883;
  assign _GEN_9082 = 11'h374 == _T_12323 ? _GEN_4 : mem_884;
  assign _GEN_9083 = 11'h375 == _T_12323 ? _GEN_4 : mem_885;
  assign _GEN_9084 = 11'h376 == _T_12323 ? _GEN_4 : mem_886;
  assign _GEN_9085 = 11'h377 == _T_12323 ? _GEN_4 : mem_887;
  assign _GEN_9086 = 11'h378 == _T_12323 ? _GEN_4 : mem_888;
  assign _GEN_9087 = 11'h379 == _T_12323 ? _GEN_4 : mem_889;
  assign _GEN_9088 = 11'h37a == _T_12323 ? _GEN_4 : mem_890;
  assign _GEN_9089 = 11'h37b == _T_12323 ? _GEN_4 : mem_891;
  assign _GEN_9090 = 11'h37c == _T_12323 ? _GEN_4 : mem_892;
  assign _GEN_9091 = 11'h37d == _T_12323 ? _GEN_4 : mem_893;
  assign _GEN_9092 = 11'h37e == _T_12323 ? _GEN_4 : mem_894;
  assign _GEN_9093 = 11'h37f == _T_12323 ? _GEN_4 : mem_895;
  assign _GEN_9094 = 11'h380 == _T_12323 ? _GEN_4 : mem_896;
  assign _GEN_9095 = 11'h381 == _T_12323 ? _GEN_4 : mem_897;
  assign _GEN_9096 = 11'h382 == _T_12323 ? _GEN_4 : mem_898;
  assign _GEN_9097 = 11'h383 == _T_12323 ? _GEN_4 : mem_899;
  assign _GEN_9098 = 11'h384 == _T_12323 ? _GEN_4 : mem_900;
  assign _GEN_9099 = 11'h385 == _T_12323 ? _GEN_4 : mem_901;
  assign _GEN_9100 = 11'h386 == _T_12323 ? _GEN_4 : mem_902;
  assign _GEN_9101 = 11'h387 == _T_12323 ? _GEN_4 : mem_903;
  assign _GEN_9102 = 11'h388 == _T_12323 ? _GEN_4 : mem_904;
  assign _GEN_9103 = 11'h389 == _T_12323 ? _GEN_4 : mem_905;
  assign _GEN_9104 = 11'h38a == _T_12323 ? _GEN_4 : mem_906;
  assign _GEN_9105 = 11'h38b == _T_12323 ? _GEN_4 : mem_907;
  assign _GEN_9106 = 11'h38c == _T_12323 ? _GEN_4 : mem_908;
  assign _GEN_9107 = 11'h38d == _T_12323 ? _GEN_4 : mem_909;
  assign _GEN_9108 = 11'h38e == _T_12323 ? _GEN_4 : mem_910;
  assign _GEN_9109 = 11'h38f == _T_12323 ? _GEN_4 : mem_911;
  assign _GEN_9110 = 11'h390 == _T_12323 ? _GEN_4 : mem_912;
  assign _GEN_9111 = 11'h391 == _T_12323 ? _GEN_4 : mem_913;
  assign _GEN_9112 = 11'h392 == _T_12323 ? _GEN_4 : mem_914;
  assign _GEN_9113 = 11'h393 == _T_12323 ? _GEN_4 : mem_915;
  assign _GEN_9114 = 11'h394 == _T_12323 ? _GEN_4 : mem_916;
  assign _GEN_9115 = 11'h395 == _T_12323 ? _GEN_4 : mem_917;
  assign _GEN_9116 = 11'h396 == _T_12323 ? _GEN_4 : mem_918;
  assign _GEN_9117 = 11'h397 == _T_12323 ? _GEN_4 : mem_919;
  assign _GEN_9118 = 11'h398 == _T_12323 ? _GEN_4 : mem_920;
  assign _GEN_9119 = 11'h399 == _T_12323 ? _GEN_4 : mem_921;
  assign _GEN_9120 = 11'h39a == _T_12323 ? _GEN_4 : mem_922;
  assign _GEN_9121 = 11'h39b == _T_12323 ? _GEN_4 : mem_923;
  assign _GEN_9122 = 11'h39c == _T_12323 ? _GEN_4 : mem_924;
  assign _GEN_9123 = 11'h39d == _T_12323 ? _GEN_4 : mem_925;
  assign _GEN_9124 = 11'h39e == _T_12323 ? _GEN_4 : mem_926;
  assign _GEN_9125 = 11'h39f == _T_12323 ? _GEN_4 : mem_927;
  assign _GEN_9126 = 11'h3a0 == _T_12323 ? _GEN_4 : mem_928;
  assign _GEN_9127 = 11'h3a1 == _T_12323 ? _GEN_4 : mem_929;
  assign _GEN_9128 = 11'h3a2 == _T_12323 ? _GEN_4 : mem_930;
  assign _GEN_9129 = 11'h3a3 == _T_12323 ? _GEN_4 : mem_931;
  assign _GEN_9130 = 11'h3a4 == _T_12323 ? _GEN_4 : mem_932;
  assign _GEN_9131 = 11'h3a5 == _T_12323 ? _GEN_4 : mem_933;
  assign _GEN_9132 = 11'h3a6 == _T_12323 ? _GEN_4 : mem_934;
  assign _GEN_9133 = 11'h3a7 == _T_12323 ? _GEN_4 : mem_935;
  assign _GEN_9134 = 11'h3a8 == _T_12323 ? _GEN_4 : mem_936;
  assign _GEN_9135 = 11'h3a9 == _T_12323 ? _GEN_4 : mem_937;
  assign _GEN_9136 = 11'h3aa == _T_12323 ? _GEN_4 : mem_938;
  assign _GEN_9137 = 11'h3ab == _T_12323 ? _GEN_4 : mem_939;
  assign _GEN_9138 = 11'h3ac == _T_12323 ? _GEN_4 : mem_940;
  assign _GEN_9139 = 11'h3ad == _T_12323 ? _GEN_4 : mem_941;
  assign _GEN_9140 = 11'h3ae == _T_12323 ? _GEN_4 : mem_942;
  assign _GEN_9141 = 11'h3af == _T_12323 ? _GEN_4 : mem_943;
  assign _GEN_9142 = 11'h3b0 == _T_12323 ? _GEN_4 : mem_944;
  assign _GEN_9143 = 11'h3b1 == _T_12323 ? _GEN_4 : mem_945;
  assign _GEN_9144 = 11'h3b2 == _T_12323 ? _GEN_4 : mem_946;
  assign _GEN_9145 = 11'h3b3 == _T_12323 ? _GEN_4 : mem_947;
  assign _GEN_9146 = 11'h3b4 == _T_12323 ? _GEN_4 : mem_948;
  assign _GEN_9147 = 11'h3b5 == _T_12323 ? _GEN_4 : mem_949;
  assign _GEN_9148 = 11'h3b6 == _T_12323 ? _GEN_4 : mem_950;
  assign _GEN_9149 = 11'h3b7 == _T_12323 ? _GEN_4 : mem_951;
  assign _GEN_9150 = 11'h3b8 == _T_12323 ? _GEN_4 : mem_952;
  assign _GEN_9151 = 11'h3b9 == _T_12323 ? _GEN_4 : mem_953;
  assign _GEN_9152 = 11'h3ba == _T_12323 ? _GEN_4 : mem_954;
  assign _GEN_9153 = 11'h3bb == _T_12323 ? _GEN_4 : mem_955;
  assign _GEN_9154 = 11'h3bc == _T_12323 ? _GEN_4 : mem_956;
  assign _GEN_9155 = 11'h3bd == _T_12323 ? _GEN_4 : mem_957;
  assign _GEN_9156 = 11'h3be == _T_12323 ? _GEN_4 : mem_958;
  assign _GEN_9157 = 11'h3bf == _T_12323 ? _GEN_4 : mem_959;
  assign _GEN_9158 = 11'h3c0 == _T_12323 ? _GEN_4 : mem_960;
  assign _GEN_9159 = 11'h3c1 == _T_12323 ? _GEN_4 : mem_961;
  assign _GEN_9160 = 11'h3c2 == _T_12323 ? _GEN_4 : mem_962;
  assign _GEN_9161 = 11'h3c3 == _T_12323 ? _GEN_4 : mem_963;
  assign _GEN_9162 = 11'h3c4 == _T_12323 ? _GEN_4 : mem_964;
  assign _GEN_9163 = 11'h3c5 == _T_12323 ? _GEN_4 : mem_965;
  assign _GEN_9164 = 11'h3c6 == _T_12323 ? _GEN_4 : mem_966;
  assign _GEN_9165 = 11'h3c7 == _T_12323 ? _GEN_4 : mem_967;
  assign _GEN_9166 = 11'h3c8 == _T_12323 ? _GEN_4 : mem_968;
  assign _GEN_9167 = 11'h3c9 == _T_12323 ? _GEN_4 : mem_969;
  assign _GEN_9168 = 11'h3ca == _T_12323 ? _GEN_4 : mem_970;
  assign _GEN_9169 = 11'h3cb == _T_12323 ? _GEN_4 : mem_971;
  assign _GEN_9170 = 11'h3cc == _T_12323 ? _GEN_4 : mem_972;
  assign _GEN_9171 = 11'h3cd == _T_12323 ? _GEN_4 : mem_973;
  assign _GEN_9172 = 11'h3ce == _T_12323 ? _GEN_4 : mem_974;
  assign _GEN_9173 = 11'h3cf == _T_12323 ? _GEN_4 : mem_975;
  assign _GEN_9174 = 11'h3d0 == _T_12323 ? _GEN_4 : mem_976;
  assign _GEN_9175 = 11'h3d1 == _T_12323 ? _GEN_4 : mem_977;
  assign _GEN_9176 = 11'h3d2 == _T_12323 ? _GEN_4 : mem_978;
  assign _GEN_9177 = 11'h3d3 == _T_12323 ? _GEN_4 : mem_979;
  assign _GEN_9178 = 11'h3d4 == _T_12323 ? _GEN_4 : mem_980;
  assign _GEN_9179 = 11'h3d5 == _T_12323 ? _GEN_4 : mem_981;
  assign _GEN_9180 = 11'h3d6 == _T_12323 ? _GEN_4 : mem_982;
  assign _GEN_9181 = 11'h3d7 == _T_12323 ? _GEN_4 : mem_983;
  assign _GEN_9182 = 11'h3d8 == _T_12323 ? _GEN_4 : mem_984;
  assign _GEN_9183 = 11'h3d9 == _T_12323 ? _GEN_4 : mem_985;
  assign _GEN_9184 = 11'h3da == _T_12323 ? _GEN_4 : mem_986;
  assign _GEN_9185 = 11'h3db == _T_12323 ? _GEN_4 : mem_987;
  assign _GEN_9186 = 11'h3dc == _T_12323 ? _GEN_4 : mem_988;
  assign _GEN_9187 = 11'h3dd == _T_12323 ? _GEN_4 : mem_989;
  assign _GEN_9188 = 11'h3de == _T_12323 ? _GEN_4 : mem_990;
  assign _GEN_9189 = 11'h3df == _T_12323 ? _GEN_4 : mem_991;
  assign _GEN_9190 = 11'h3e0 == _T_12323 ? _GEN_4 : mem_992;
  assign _GEN_9191 = 11'h3e1 == _T_12323 ? _GEN_4 : mem_993;
  assign _GEN_9192 = 11'h3e2 == _T_12323 ? _GEN_4 : mem_994;
  assign _GEN_9193 = 11'h3e3 == _T_12323 ? _GEN_4 : mem_995;
  assign _GEN_9194 = 11'h3e4 == _T_12323 ? _GEN_4 : mem_996;
  assign _GEN_9195 = 11'h3e5 == _T_12323 ? _GEN_4 : mem_997;
  assign _GEN_9196 = 11'h3e6 == _T_12323 ? _GEN_4 : mem_998;
  assign _GEN_9197 = 11'h3e7 == _T_12323 ? _GEN_4 : mem_999;
  assign _GEN_9198 = 11'h3e8 == _T_12323 ? _GEN_4 : mem_1000;
  assign _GEN_9199 = 11'h3e9 == _T_12323 ? _GEN_4 : mem_1001;
  assign _GEN_9200 = 11'h3ea == _T_12323 ? _GEN_4 : mem_1002;
  assign _GEN_9201 = 11'h3eb == _T_12323 ? _GEN_4 : mem_1003;
  assign _GEN_9202 = 11'h3ec == _T_12323 ? _GEN_4 : mem_1004;
  assign _GEN_9203 = 11'h3ed == _T_12323 ? _GEN_4 : mem_1005;
  assign _GEN_9204 = 11'h3ee == _T_12323 ? _GEN_4 : mem_1006;
  assign _GEN_9205 = 11'h3ef == _T_12323 ? _GEN_4 : mem_1007;
  assign _GEN_9206 = 11'h3f0 == _T_12323 ? _GEN_4 : mem_1008;
  assign _GEN_9207 = 11'h3f1 == _T_12323 ? _GEN_4 : mem_1009;
  assign _GEN_9208 = 11'h3f2 == _T_12323 ? _GEN_4 : mem_1010;
  assign _GEN_9209 = 11'h3f3 == _T_12323 ? _GEN_4 : mem_1011;
  assign _GEN_9210 = 11'h3f4 == _T_12323 ? _GEN_4 : mem_1012;
  assign _GEN_9211 = 11'h3f5 == _T_12323 ? _GEN_4 : mem_1013;
  assign _GEN_9212 = 11'h3f6 == _T_12323 ? _GEN_4 : mem_1014;
  assign _GEN_9213 = 11'h3f7 == _T_12323 ? _GEN_4 : mem_1015;
  assign _GEN_9214 = 11'h3f8 == _T_12323 ? _GEN_4 : mem_1016;
  assign _GEN_9215 = 11'h3f9 == _T_12323 ? _GEN_4 : mem_1017;
  assign _GEN_9216 = 11'h3fa == _T_12323 ? _GEN_4 : mem_1018;
  assign _GEN_9217 = 11'h3fb == _T_12323 ? _GEN_4 : mem_1019;
  assign _GEN_9218 = 11'h3fc == _T_12323 ? _GEN_4 : mem_1020;
  assign _GEN_9219 = 11'h3fd == _T_12323 ? _GEN_4 : mem_1021;
  assign _GEN_9220 = 11'h3fe == _T_12323 ? _GEN_4 : mem_1022;
  assign _GEN_9221 = 11'h3ff == _T_12323 ? _GEN_4 : mem_1023;
  assign _GEN_9222 = 11'h400 == _T_12323 ? _GEN_4 : mem_1024;
  assign _GEN_9223 = 11'h401 == _T_12323 ? _GEN_4 : mem_1025;
  assign _GEN_9224 = 11'h402 == _T_12323 ? _GEN_4 : mem_1026;
  assign _GEN_9225 = 11'h403 == _T_12323 ? _GEN_4 : mem_1027;
  assign _GEN_9226 = 11'h404 == _T_12323 ? _GEN_4 : mem_1028;
  assign _GEN_9227 = 11'h405 == _T_12323 ? _GEN_4 : mem_1029;
  assign _GEN_9228 = 11'h406 == _T_12323 ? _GEN_4 : mem_1030;
  assign _GEN_9229 = 11'h407 == _T_12323 ? _GEN_4 : mem_1031;
  assign _GEN_9230 = 11'h408 == _T_12323 ? _GEN_4 : mem_1032;
  assign _GEN_9231 = 11'h409 == _T_12323 ? _GEN_4 : mem_1033;
  assign _GEN_9232 = 11'h40a == _T_12323 ? _GEN_4 : mem_1034;
  assign _GEN_9233 = 11'h40b == _T_12323 ? _GEN_4 : mem_1035;
  assign _GEN_9234 = 11'h40c == _T_12323 ? _GEN_4 : mem_1036;
  assign _GEN_9235 = 11'h40d == _T_12323 ? _GEN_4 : mem_1037;
  assign _GEN_9236 = 11'h40e == _T_12323 ? _GEN_4 : mem_1038;
  assign _GEN_9237 = 11'h40f == _T_12323 ? _GEN_4 : mem_1039;
  assign _GEN_9238 = 11'h410 == _T_12323 ? _GEN_4 : mem_1040;
  assign _GEN_9239 = 11'h411 == _T_12323 ? _GEN_4 : mem_1041;
  assign _GEN_9240 = 11'h412 == _T_12323 ? _GEN_4 : mem_1042;
  assign _GEN_9241 = 11'h413 == _T_12323 ? _GEN_4 : mem_1043;
  assign _GEN_9242 = 11'h414 == _T_12323 ? _GEN_4 : mem_1044;
  assign _GEN_9243 = 11'h415 == _T_12323 ? _GEN_4 : mem_1045;
  assign _GEN_9244 = 11'h416 == _T_12323 ? _GEN_4 : mem_1046;
  assign _GEN_9245 = 11'h417 == _T_12323 ? _GEN_4 : mem_1047;
  assign _GEN_9246 = 11'h418 == _T_12323 ? _GEN_4 : mem_1048;
  assign _GEN_9247 = 11'h419 == _T_12323 ? _GEN_4 : mem_1049;
  assign _GEN_9248 = 11'h41a == _T_12323 ? _GEN_4 : mem_1050;
  assign _GEN_9249 = 11'h41b == _T_12323 ? _GEN_4 : mem_1051;
  assign _GEN_9250 = 11'h41c == _T_12323 ? _GEN_4 : mem_1052;
  assign _GEN_9251 = 11'h41d == _T_12323 ? _GEN_4 : mem_1053;
  assign _GEN_9252 = 11'h41e == _T_12323 ? _GEN_4 : mem_1054;
  assign _GEN_9253 = 11'h41f == _T_12323 ? _GEN_4 : mem_1055;
  assign _GEN_9254 = 11'h420 == _T_12323 ? _GEN_4 : mem_1056;
  assign _GEN_9255 = 11'h421 == _T_12323 ? _GEN_4 : mem_1057;
  assign _GEN_9256 = 11'h422 == _T_12323 ? _GEN_4 : mem_1058;
  assign _GEN_9257 = 11'h423 == _T_12323 ? _GEN_4 : mem_1059;
  assign _GEN_9258 = 11'h424 == _T_12323 ? _GEN_4 : mem_1060;
  assign _GEN_9259 = 11'h425 == _T_12323 ? _GEN_4 : mem_1061;
  assign _GEN_9260 = 11'h426 == _T_12323 ? _GEN_4 : mem_1062;
  assign _GEN_9261 = 11'h427 == _T_12323 ? _GEN_4 : mem_1063;
  assign _GEN_9262 = 11'h428 == _T_12323 ? _GEN_4 : mem_1064;
  assign _GEN_9263 = 11'h429 == _T_12323 ? _GEN_4 : mem_1065;
  assign _GEN_9264 = 11'h42a == _T_12323 ? _GEN_4 : mem_1066;
  assign _GEN_9265 = 11'h42b == _T_12323 ? _GEN_4 : mem_1067;
  assign _GEN_9266 = 11'h42c == _T_12323 ? _GEN_4 : mem_1068;
  assign _GEN_9267 = 11'h42d == _T_12323 ? _GEN_4 : mem_1069;
  assign _GEN_9268 = 11'h42e == _T_12323 ? _GEN_4 : mem_1070;
  assign _GEN_9269 = 11'h42f == _T_12323 ? _GEN_4 : mem_1071;
  assign _GEN_9270 = 11'h430 == _T_12323 ? _GEN_4 : mem_1072;
  assign _GEN_9271 = 11'h431 == _T_12323 ? _GEN_4 : mem_1073;
  assign _GEN_9272 = 11'h432 == _T_12323 ? _GEN_4 : mem_1074;
  assign _GEN_9273 = 11'h433 == _T_12323 ? _GEN_4 : mem_1075;
  assign _GEN_9274 = 11'h434 == _T_12323 ? _GEN_4 : mem_1076;
  assign _GEN_9275 = 11'h435 == _T_12323 ? _GEN_4 : mem_1077;
  assign _GEN_9276 = 11'h436 == _T_12323 ? _GEN_4 : mem_1078;
  assign _GEN_9277 = 11'h437 == _T_12323 ? _GEN_4 : mem_1079;
  assign _GEN_9278 = 11'h438 == _T_12323 ? _GEN_4 : mem_1080;
  assign _GEN_9279 = 11'h439 == _T_12323 ? _GEN_4 : mem_1081;
  assign _GEN_9280 = 11'h43a == _T_12323 ? _GEN_4 : mem_1082;
  assign _GEN_9281 = 11'h43b == _T_12323 ? _GEN_4 : mem_1083;
  assign _GEN_9282 = 11'h43c == _T_12323 ? _GEN_4 : mem_1084;
  assign _GEN_9283 = 11'h43d == _T_12323 ? _GEN_4 : mem_1085;
  assign _GEN_9284 = 11'h43e == _T_12323 ? _GEN_4 : mem_1086;
  assign _GEN_9285 = 11'h43f == _T_12323 ? _GEN_4 : mem_1087;
  assign _GEN_9286 = 11'h440 == _T_12323 ? _GEN_4 : mem_1088;
  assign _GEN_9287 = 11'h441 == _T_12323 ? _GEN_4 : mem_1089;
  assign _GEN_9288 = 11'h442 == _T_12323 ? _GEN_4 : mem_1090;
  assign _GEN_9289 = 11'h443 == _T_12323 ? _GEN_4 : mem_1091;
  assign _GEN_9290 = 11'h444 == _T_12323 ? _GEN_4 : mem_1092;
  assign _GEN_9291 = 11'h445 == _T_12323 ? _GEN_4 : mem_1093;
  assign _GEN_9292 = 11'h446 == _T_12323 ? _GEN_4 : mem_1094;
  assign _GEN_9293 = 11'h447 == _T_12323 ? _GEN_4 : mem_1095;
  assign _GEN_9294 = 11'h448 == _T_12323 ? _GEN_4 : mem_1096;
  assign _GEN_9295 = 11'h449 == _T_12323 ? _GEN_4 : mem_1097;
  assign _GEN_9296 = 11'h44a == _T_12323 ? _GEN_4 : mem_1098;
  assign _GEN_9297 = 11'h44b == _T_12323 ? _GEN_4 : mem_1099;
  assign _GEN_9298 = 11'h44c == _T_12323 ? _GEN_4 : mem_1100;
  assign _GEN_9299 = 11'h44d == _T_12323 ? _GEN_4 : mem_1101;
  assign _GEN_9300 = 11'h44e == _T_12323 ? _GEN_4 : mem_1102;
  assign _GEN_9301 = 11'h44f == _T_12323 ? _GEN_4 : mem_1103;
  assign _GEN_9302 = 11'h450 == _T_12323 ? _GEN_4 : mem_1104;
  assign _GEN_9303 = 11'h451 == _T_12323 ? _GEN_4 : mem_1105;
  assign _GEN_9304 = 11'h452 == _T_12323 ? _GEN_4 : mem_1106;
  assign _GEN_9305 = 11'h453 == _T_12323 ? _GEN_4 : mem_1107;
  assign _GEN_9306 = 11'h454 == _T_12323 ? _GEN_4 : mem_1108;
  assign _GEN_9307 = 11'h455 == _T_12323 ? _GEN_4 : mem_1109;
  assign _GEN_9308 = 11'h456 == _T_12323 ? _GEN_4 : mem_1110;
  assign _GEN_9309 = 11'h457 == _T_12323 ? _GEN_4 : mem_1111;
  assign _GEN_9310 = 11'h458 == _T_12323 ? _GEN_4 : mem_1112;
  assign _GEN_9311 = 11'h459 == _T_12323 ? _GEN_4 : mem_1113;
  assign _GEN_9312 = 11'h45a == _T_12323 ? _GEN_4 : mem_1114;
  assign _GEN_9313 = 11'h45b == _T_12323 ? _GEN_4 : mem_1115;
  assign _GEN_9314 = 11'h45c == _T_12323 ? _GEN_4 : mem_1116;
  assign _GEN_9315 = 11'h45d == _T_12323 ? _GEN_4 : mem_1117;
  assign _GEN_9316 = 11'h45e == _T_12323 ? _GEN_4 : mem_1118;
  assign _GEN_9317 = 11'h45f == _T_12323 ? _GEN_4 : mem_1119;
  assign _GEN_9318 = 11'h460 == _T_12323 ? _GEN_4 : mem_1120;
  assign _GEN_9319 = 11'h461 == _T_12323 ? _GEN_4 : mem_1121;
  assign _GEN_9320 = 11'h462 == _T_12323 ? _GEN_4 : mem_1122;
  assign _GEN_9321 = 11'h463 == _T_12323 ? _GEN_4 : mem_1123;
  assign _GEN_9322 = 11'h464 == _T_12323 ? _GEN_4 : mem_1124;
  assign _GEN_9323 = 11'h465 == _T_12323 ? _GEN_4 : mem_1125;
  assign _GEN_9324 = 11'h466 == _T_12323 ? _GEN_4 : mem_1126;
  assign _GEN_9325 = 11'h467 == _T_12323 ? _GEN_4 : mem_1127;
  assign _GEN_9326 = 11'h468 == _T_12323 ? _GEN_4 : mem_1128;
  assign _GEN_9327 = 11'h469 == _T_12323 ? _GEN_4 : mem_1129;
  assign _GEN_9328 = 11'h46a == _T_12323 ? _GEN_4 : mem_1130;
  assign _GEN_9329 = 11'h46b == _T_12323 ? _GEN_4 : mem_1131;
  assign _GEN_9330 = 11'h46c == _T_12323 ? _GEN_4 : mem_1132;
  assign _GEN_9331 = 11'h46d == _T_12323 ? _GEN_4 : mem_1133;
  assign _GEN_9332 = 11'h46e == _T_12323 ? _GEN_4 : mem_1134;
  assign _GEN_9333 = 11'h46f == _T_12323 ? _GEN_4 : mem_1135;
  assign _GEN_9334 = 11'h470 == _T_12323 ? _GEN_4 : mem_1136;
  assign _GEN_9335 = 11'h471 == _T_12323 ? _GEN_4 : mem_1137;
  assign _GEN_9336 = 11'h472 == _T_12323 ? _GEN_4 : mem_1138;
  assign _GEN_9337 = 11'h473 == _T_12323 ? _GEN_4 : mem_1139;
  assign _GEN_9338 = 11'h474 == _T_12323 ? _GEN_4 : mem_1140;
  assign _GEN_9339 = 11'h475 == _T_12323 ? _GEN_4 : mem_1141;
  assign _GEN_9340 = 11'h476 == _T_12323 ? _GEN_4 : mem_1142;
  assign _GEN_9341 = 11'h477 == _T_12323 ? _GEN_4 : mem_1143;
  assign _GEN_9342 = 11'h478 == _T_12323 ? _GEN_4 : mem_1144;
  assign _GEN_9343 = 11'h479 == _T_12323 ? _GEN_4 : mem_1145;
  assign _GEN_9344 = 11'h47a == _T_12323 ? _GEN_4 : mem_1146;
  assign _GEN_9345 = 11'h47b == _T_12323 ? _GEN_4 : mem_1147;
  assign _GEN_9346 = 11'h47c == _T_12323 ? _GEN_4 : mem_1148;
  assign _GEN_9347 = 11'h47d == _T_12323 ? _GEN_4 : mem_1149;
  assign _GEN_9348 = 11'h47e == _T_12323 ? _GEN_4 : mem_1150;
  assign _GEN_9349 = 11'h47f == _T_12323 ? _GEN_4 : mem_1151;
  assign _GEN_9350 = 11'h480 == _T_12323 ? _GEN_4 : mem_1152;
  assign _GEN_9351 = 11'h481 == _T_12323 ? _GEN_4 : mem_1153;
  assign _GEN_9352 = 11'h482 == _T_12323 ? _GEN_4 : mem_1154;
  assign _GEN_9353 = 11'h483 == _T_12323 ? _GEN_4 : mem_1155;
  assign _GEN_9354 = 11'h484 == _T_12323 ? _GEN_4 : mem_1156;
  assign _GEN_9355 = 11'h485 == _T_12323 ? _GEN_4 : mem_1157;
  assign _GEN_9356 = 11'h486 == _T_12323 ? _GEN_4 : mem_1158;
  assign _GEN_9357 = 11'h487 == _T_12323 ? _GEN_4 : mem_1159;
  assign _GEN_9358 = 11'h488 == _T_12323 ? _GEN_4 : mem_1160;
  assign _GEN_9359 = 11'h489 == _T_12323 ? _GEN_4 : mem_1161;
  assign _GEN_9360 = 11'h48a == _T_12323 ? _GEN_4 : mem_1162;
  assign _GEN_9361 = 11'h48b == _T_12323 ? _GEN_4 : mem_1163;
  assign _GEN_9362 = 11'h48c == _T_12323 ? _GEN_4 : mem_1164;
  assign _GEN_9363 = 11'h48d == _T_12323 ? _GEN_4 : mem_1165;
  assign _GEN_9364 = 11'h48e == _T_12323 ? _GEN_4 : mem_1166;
  assign _GEN_9365 = 11'h48f == _T_12323 ? _GEN_4 : mem_1167;
  assign _GEN_9366 = 11'h490 == _T_12323 ? _GEN_4 : mem_1168;
  assign _GEN_9367 = 11'h491 == _T_12323 ? _GEN_4 : mem_1169;
  assign _GEN_9368 = 11'h492 == _T_12323 ? _GEN_4 : mem_1170;
  assign _GEN_9369 = 11'h493 == _T_12323 ? _GEN_4 : mem_1171;
  assign _GEN_9370 = 11'h494 == _T_12323 ? _GEN_4 : mem_1172;
  assign _GEN_9371 = 11'h495 == _T_12323 ? _GEN_4 : mem_1173;
  assign _GEN_9372 = 11'h496 == _T_12323 ? _GEN_4 : mem_1174;
  assign _GEN_9373 = 11'h497 == _T_12323 ? _GEN_4 : mem_1175;
  assign _GEN_9374 = 11'h498 == _T_12323 ? _GEN_4 : mem_1176;
  assign _GEN_9375 = 11'h499 == _T_12323 ? _GEN_4 : mem_1177;
  assign _GEN_9376 = 11'h49a == _T_12323 ? _GEN_4 : mem_1178;
  assign _GEN_9377 = 11'h49b == _T_12323 ? _GEN_4 : mem_1179;
  assign _GEN_9378 = 11'h49c == _T_12323 ? _GEN_4 : mem_1180;
  assign _GEN_9379 = 11'h49d == _T_12323 ? _GEN_4 : mem_1181;
  assign _GEN_9380 = 11'h49e == _T_12323 ? _GEN_4 : mem_1182;
  assign _GEN_9381 = 11'h49f == _T_12323 ? _GEN_4 : mem_1183;
  assign _GEN_9382 = 11'h4a0 == _T_12323 ? _GEN_4 : mem_1184;
  assign _GEN_9383 = 11'h4a1 == _T_12323 ? _GEN_4 : mem_1185;
  assign _GEN_9384 = 11'h4a2 == _T_12323 ? _GEN_4 : mem_1186;
  assign _GEN_9385 = 11'h4a3 == _T_12323 ? _GEN_4 : mem_1187;
  assign _GEN_9386 = 11'h4a4 == _T_12323 ? _GEN_4 : mem_1188;
  assign _GEN_9387 = 11'h4a5 == _T_12323 ? _GEN_4 : mem_1189;
  assign _GEN_9388 = 11'h4a6 == _T_12323 ? _GEN_4 : mem_1190;
  assign _GEN_9389 = 11'h4a7 == _T_12323 ? _GEN_4 : mem_1191;
  assign _GEN_9390 = 11'h4a8 == _T_12323 ? _GEN_4 : mem_1192;
  assign _GEN_9391 = 11'h4a9 == _T_12323 ? _GEN_4 : mem_1193;
  assign _GEN_9392 = 11'h4aa == _T_12323 ? _GEN_4 : mem_1194;
  assign _GEN_9393 = 11'h4ab == _T_12323 ? _GEN_4 : mem_1195;
  assign _GEN_9394 = 11'h4ac == _T_12323 ? _GEN_4 : mem_1196;
  assign _GEN_9395 = 11'h4ad == _T_12323 ? _GEN_4 : mem_1197;
  assign _GEN_9396 = 11'h4ae == _T_12323 ? _GEN_4 : mem_1198;
  assign _GEN_9397 = 11'h4af == _T_12323 ? _GEN_4 : mem_1199;
  assign _GEN_9398 = 11'h4b0 == _T_12323 ? _GEN_4 : mem_1200;
  assign _GEN_9399 = 11'h4b1 == _T_12323 ? _GEN_4 : mem_1201;
  assign _GEN_9400 = 11'h4b2 == _T_12323 ? _GEN_4 : mem_1202;
  assign _GEN_9401 = 11'h4b3 == _T_12323 ? _GEN_4 : mem_1203;
  assign _GEN_9402 = 11'h4b4 == _T_12323 ? _GEN_4 : mem_1204;
  assign _GEN_9403 = 11'h4b5 == _T_12323 ? _GEN_4 : mem_1205;
  assign _GEN_9404 = 11'h4b6 == _T_12323 ? _GEN_4 : mem_1206;
  assign _GEN_9405 = 11'h4b7 == _T_12323 ? _GEN_4 : mem_1207;
  assign _GEN_9406 = 11'h4b8 == _T_12323 ? _GEN_4 : mem_1208;
  assign _GEN_9407 = 11'h4b9 == _T_12323 ? _GEN_4 : mem_1209;
  assign _GEN_9408 = 11'h4ba == _T_12323 ? _GEN_4 : mem_1210;
  assign _GEN_9409 = 11'h4bb == _T_12323 ? _GEN_4 : mem_1211;
  assign _GEN_9410 = 11'h4bc == _T_12323 ? _GEN_4 : mem_1212;
  assign _GEN_9411 = 11'h4bd == _T_12323 ? _GEN_4 : mem_1213;
  assign _GEN_9412 = 11'h4be == _T_12323 ? _GEN_4 : mem_1214;
  assign _GEN_9413 = 11'h4bf == _T_12323 ? _GEN_4 : mem_1215;
  assign _GEN_9414 = 11'h4c0 == _T_12323 ? _GEN_4 : mem_1216;
  assign _GEN_9415 = 11'h4c1 == _T_12323 ? _GEN_4 : mem_1217;
  assign _GEN_9416 = 11'h4c2 == _T_12323 ? _GEN_4 : mem_1218;
  assign _GEN_9417 = 11'h4c3 == _T_12323 ? _GEN_4 : mem_1219;
  assign _GEN_9418 = 11'h4c4 == _T_12323 ? _GEN_4 : mem_1220;
  assign _GEN_9419 = 11'h4c5 == _T_12323 ? _GEN_4 : mem_1221;
  assign _GEN_9420 = 11'h4c6 == _T_12323 ? _GEN_4 : mem_1222;
  assign _GEN_9421 = 11'h4c7 == _T_12323 ? _GEN_4 : mem_1223;
  assign _GEN_9422 = 11'h4c8 == _T_12323 ? _GEN_4 : mem_1224;
  assign _GEN_9423 = 11'h4c9 == _T_12323 ? _GEN_4 : mem_1225;
  assign _GEN_9424 = 11'h4ca == _T_12323 ? _GEN_4 : mem_1226;
  assign _GEN_9425 = 11'h4cb == _T_12323 ? _GEN_4 : mem_1227;
  assign _GEN_9426 = 11'h4cc == _T_12323 ? _GEN_4 : mem_1228;
  assign _GEN_9427 = 11'h4cd == _T_12323 ? _GEN_4 : mem_1229;
  assign _GEN_9428 = 11'h4ce == _T_12323 ? _GEN_4 : mem_1230;
  assign _GEN_9429 = 11'h4cf == _T_12323 ? _GEN_4 : mem_1231;
  assign _GEN_9430 = 11'h4d0 == _T_12323 ? _GEN_4 : mem_1232;
  assign _GEN_9431 = 11'h4d1 == _T_12323 ? _GEN_4 : mem_1233;
  assign _GEN_9432 = 11'h4d2 == _T_12323 ? _GEN_4 : mem_1234;
  assign _GEN_9433 = 11'h4d3 == _T_12323 ? _GEN_4 : mem_1235;
  assign _GEN_9434 = 11'h4d4 == _T_12323 ? _GEN_4 : mem_1236;
  assign _GEN_9435 = 11'h4d5 == _T_12323 ? _GEN_4 : mem_1237;
  assign _GEN_9436 = 11'h4d6 == _T_12323 ? _GEN_4 : mem_1238;
  assign _GEN_9437 = 11'h4d7 == _T_12323 ? _GEN_4 : mem_1239;
  assign _GEN_9438 = 11'h4d8 == _T_12323 ? _GEN_4 : mem_1240;
  assign _GEN_9439 = 11'h4d9 == _T_12323 ? _GEN_4 : mem_1241;
  assign _GEN_9440 = 11'h4da == _T_12323 ? _GEN_4 : mem_1242;
  assign _GEN_9441 = 11'h4db == _T_12323 ? _GEN_4 : mem_1243;
  assign _GEN_9442 = 11'h4dc == _T_12323 ? _GEN_4 : mem_1244;
  assign _GEN_9443 = 11'h4dd == _T_12323 ? _GEN_4 : mem_1245;
  assign _GEN_9444 = 11'h4de == _T_12323 ? _GEN_4 : mem_1246;
  assign _GEN_9445 = 11'h4df == _T_12323 ? _GEN_4 : mem_1247;
  assign _GEN_9446 = 11'h4e0 == _T_12323 ? _GEN_4 : mem_1248;
  assign _GEN_9447 = 11'h4e1 == _T_12323 ? _GEN_4 : mem_1249;
  assign _GEN_9448 = 11'h4e2 == _T_12323 ? _GEN_4 : mem_1250;
  assign _GEN_9449 = 11'h4e3 == _T_12323 ? _GEN_4 : mem_1251;
  assign _GEN_9450 = 11'h4e4 == _T_12323 ? _GEN_4 : mem_1252;
  assign _GEN_9451 = 11'h4e5 == _T_12323 ? _GEN_4 : mem_1253;
  assign _GEN_9452 = 11'h4e6 == _T_12323 ? _GEN_4 : mem_1254;
  assign _GEN_9453 = 11'h4e7 == _T_12323 ? _GEN_4 : mem_1255;
  assign _GEN_9454 = 11'h4e8 == _T_12323 ? _GEN_4 : mem_1256;
  assign _GEN_9455 = 11'h4e9 == _T_12323 ? _GEN_4 : mem_1257;
  assign _GEN_9456 = 11'h4ea == _T_12323 ? _GEN_4 : mem_1258;
  assign _GEN_9457 = 11'h4eb == _T_12323 ? _GEN_4 : mem_1259;
  assign _GEN_9458 = 11'h4ec == _T_12323 ? _GEN_4 : mem_1260;
  assign _GEN_9459 = 11'h4ed == _T_12323 ? _GEN_4 : mem_1261;
  assign _GEN_9460 = 11'h4ee == _T_12323 ? _GEN_4 : mem_1262;
  assign _GEN_9461 = 11'h4ef == _T_12323 ? _GEN_4 : mem_1263;
  assign _GEN_9462 = 11'h4f0 == _T_12323 ? _GEN_4 : mem_1264;
  assign _GEN_9463 = 11'h4f1 == _T_12323 ? _GEN_4 : mem_1265;
  assign _GEN_9464 = 11'h4f2 == _T_12323 ? _GEN_4 : mem_1266;
  assign _GEN_9465 = 11'h4f3 == _T_12323 ? _GEN_4 : mem_1267;
  assign _GEN_9466 = 11'h4f4 == _T_12323 ? _GEN_4 : mem_1268;
  assign _GEN_9467 = 11'h4f5 == _T_12323 ? _GEN_4 : mem_1269;
  assign _GEN_9468 = 11'h4f6 == _T_12323 ? _GEN_4 : mem_1270;
  assign _GEN_9469 = 11'h4f7 == _T_12323 ? _GEN_4 : mem_1271;
  assign _GEN_9470 = 11'h4f8 == _T_12323 ? _GEN_4 : mem_1272;
  assign _GEN_9471 = 11'h4f9 == _T_12323 ? _GEN_4 : mem_1273;
  assign _GEN_9472 = 11'h4fa == _T_12323 ? _GEN_4 : mem_1274;
  assign _GEN_9473 = 11'h4fb == _T_12323 ? _GEN_4 : mem_1275;
  assign _GEN_9474 = 11'h4fc == _T_12323 ? _GEN_4 : mem_1276;
  assign _GEN_9475 = 11'h4fd == _T_12323 ? _GEN_4 : mem_1277;
  assign _GEN_9476 = 11'h4fe == _T_12323 ? _GEN_4 : mem_1278;
  assign _GEN_9477 = 11'h4ff == _T_12323 ? _GEN_4 : mem_1279;
  assign _GEN_9478 = 11'h500 == _T_12323 ? _GEN_4 : mem_1280;
  assign _GEN_9479 = 11'h501 == _T_12323 ? _GEN_4 : mem_1281;
  assign _GEN_9480 = 11'h502 == _T_12323 ? _GEN_4 : mem_1282;
  assign _GEN_9481 = 11'h503 == _T_12323 ? _GEN_4 : mem_1283;
  assign _GEN_9482 = 11'h504 == _T_12323 ? _GEN_4 : mem_1284;
  assign _GEN_9483 = 11'h505 == _T_12323 ? _GEN_4 : mem_1285;
  assign _GEN_9484 = 11'h506 == _T_12323 ? _GEN_4 : mem_1286;
  assign _GEN_9485 = 11'h507 == _T_12323 ? _GEN_4 : mem_1287;
  assign _GEN_9486 = 11'h508 == _T_12323 ? _GEN_4 : mem_1288;
  assign _GEN_9487 = 11'h509 == _T_12323 ? _GEN_4 : mem_1289;
  assign _GEN_9488 = 11'h50a == _T_12323 ? _GEN_4 : mem_1290;
  assign _GEN_9489 = 11'h50b == _T_12323 ? _GEN_4 : mem_1291;
  assign _GEN_9490 = 11'h50c == _T_12323 ? _GEN_4 : mem_1292;
  assign _GEN_9491 = 11'h50d == _T_12323 ? _GEN_4 : mem_1293;
  assign _GEN_9492 = 11'h50e == _T_12323 ? _GEN_4 : mem_1294;
  assign _GEN_9493 = 11'h50f == _T_12323 ? _GEN_4 : mem_1295;
  assign _GEN_9494 = 11'h510 == _T_12323 ? _GEN_4 : mem_1296;
  assign _GEN_9495 = 11'h511 == _T_12323 ? _GEN_4 : mem_1297;
  assign _GEN_9496 = 11'h512 == _T_12323 ? _GEN_4 : mem_1298;
  assign _GEN_9497 = 11'h513 == _T_12323 ? _GEN_4 : mem_1299;
  assign _GEN_9498 = 11'h514 == _T_12323 ? _GEN_4 : mem_1300;
  assign _GEN_9499 = 11'h515 == _T_12323 ? _GEN_4 : mem_1301;
  assign _GEN_9500 = 11'h516 == _T_12323 ? _GEN_4 : mem_1302;
  assign _GEN_9501 = 11'h517 == _T_12323 ? _GEN_4 : mem_1303;
  assign _GEN_9502 = 11'h518 == _T_12323 ? _GEN_4 : mem_1304;
  assign _GEN_9503 = 11'h519 == _T_12323 ? _GEN_4 : mem_1305;
  assign _GEN_9504 = 11'h51a == _T_12323 ? _GEN_4 : mem_1306;
  assign _GEN_9505 = 11'h51b == _T_12323 ? _GEN_4 : mem_1307;
  assign _GEN_9506 = 11'h51c == _T_12323 ? _GEN_4 : mem_1308;
  assign _GEN_9507 = 11'h51d == _T_12323 ? _GEN_4 : mem_1309;
  assign _GEN_9508 = 11'h51e == _T_12323 ? _GEN_4 : mem_1310;
  assign _GEN_9509 = 11'h51f == _T_12323 ? _GEN_4 : mem_1311;
  assign _GEN_9510 = 11'h520 == _T_12323 ? _GEN_4 : mem_1312;
  assign _GEN_9511 = 11'h521 == _T_12323 ? _GEN_4 : mem_1313;
  assign _GEN_9512 = 11'h522 == _T_12323 ? _GEN_4 : mem_1314;
  assign _GEN_9513 = 11'h523 == _T_12323 ? _GEN_4 : mem_1315;
  assign _GEN_9514 = 11'h524 == _T_12323 ? _GEN_4 : mem_1316;
  assign _GEN_9515 = 11'h525 == _T_12323 ? _GEN_4 : mem_1317;
  assign _GEN_9516 = 11'h526 == _T_12323 ? _GEN_4 : mem_1318;
  assign _GEN_9517 = 11'h527 == _T_12323 ? _GEN_4 : mem_1319;
  assign _GEN_9518 = 11'h528 == _T_12323 ? _GEN_4 : mem_1320;
  assign _GEN_9519 = 11'h529 == _T_12323 ? _GEN_4 : mem_1321;
  assign _GEN_9520 = 11'h52a == _T_12323 ? _GEN_4 : mem_1322;
  assign _GEN_9521 = 11'h52b == _T_12323 ? _GEN_4 : mem_1323;
  assign _GEN_9522 = 11'h52c == _T_12323 ? _GEN_4 : mem_1324;
  assign _GEN_9523 = 11'h52d == _T_12323 ? _GEN_4 : mem_1325;
  assign _GEN_9524 = 11'h52e == _T_12323 ? _GEN_4 : mem_1326;
  assign _GEN_9525 = 11'h52f == _T_12323 ? _GEN_4 : mem_1327;
  assign _GEN_9526 = 11'h530 == _T_12323 ? _GEN_4 : mem_1328;
  assign _GEN_9527 = 11'h531 == _T_12323 ? _GEN_4 : mem_1329;
  assign _GEN_9528 = 11'h532 == _T_12323 ? _GEN_4 : mem_1330;
  assign _GEN_9529 = 11'h533 == _T_12323 ? _GEN_4 : mem_1331;
  assign _GEN_9530 = 11'h534 == _T_12323 ? _GEN_4 : mem_1332;
  assign _GEN_9531 = 11'h535 == _T_12323 ? _GEN_4 : mem_1333;
  assign _GEN_9532 = 11'h536 == _T_12323 ? _GEN_4 : mem_1334;
  assign _GEN_9533 = 11'h537 == _T_12323 ? _GEN_4 : mem_1335;
  assign _GEN_9534 = 11'h538 == _T_12323 ? _GEN_4 : mem_1336;
  assign _GEN_9535 = 11'h539 == _T_12323 ? _GEN_4 : mem_1337;
  assign _GEN_9536 = 11'h53a == _T_12323 ? _GEN_4 : mem_1338;
  assign _GEN_9537 = 11'h53b == _T_12323 ? _GEN_4 : mem_1339;
  assign _GEN_9538 = 11'h53c == _T_12323 ? _GEN_4 : mem_1340;
  assign _GEN_9539 = 11'h53d == _T_12323 ? _GEN_4 : mem_1341;
  assign _GEN_9540 = 11'h53e == _T_12323 ? _GEN_4 : mem_1342;
  assign _GEN_9541 = 11'h53f == _T_12323 ? _GEN_4 : mem_1343;
  assign _GEN_9542 = 11'h540 == _T_12323 ? _GEN_4 : mem_1344;
  assign _GEN_9543 = 11'h541 == _T_12323 ? _GEN_4 : mem_1345;
  assign _GEN_9544 = 11'h542 == _T_12323 ? _GEN_4 : mem_1346;
  assign _GEN_9545 = 11'h543 == _T_12323 ? _GEN_4 : mem_1347;
  assign _GEN_9546 = 11'h544 == _T_12323 ? _GEN_4 : mem_1348;
  assign _GEN_9547 = 11'h545 == _T_12323 ? _GEN_4 : mem_1349;
  assign _GEN_9548 = 11'h546 == _T_12323 ? _GEN_4 : mem_1350;
  assign _GEN_9549 = 11'h547 == _T_12323 ? _GEN_4 : mem_1351;
  assign _GEN_9550 = 11'h548 == _T_12323 ? _GEN_4 : mem_1352;
  assign _GEN_9551 = 11'h549 == _T_12323 ? _GEN_4 : mem_1353;
  assign _GEN_9552 = 11'h54a == _T_12323 ? _GEN_4 : mem_1354;
  assign _GEN_9553 = 11'h54b == _T_12323 ? _GEN_4 : mem_1355;
  assign _GEN_9554 = 11'h54c == _T_12323 ? _GEN_4 : mem_1356;
  assign _GEN_9555 = 11'h54d == _T_12323 ? _GEN_4 : mem_1357;
  assign _GEN_9556 = 11'h54e == _T_12323 ? _GEN_4 : mem_1358;
  assign _GEN_9557 = 11'h54f == _T_12323 ? _GEN_4 : mem_1359;
  assign _GEN_9558 = 11'h550 == _T_12323 ? _GEN_4 : mem_1360;
  assign _GEN_9559 = 11'h551 == _T_12323 ? _GEN_4 : mem_1361;
  assign _GEN_9560 = 11'h552 == _T_12323 ? _GEN_4 : mem_1362;
  assign _GEN_9561 = 11'h553 == _T_12323 ? _GEN_4 : mem_1363;
  assign _GEN_9562 = 11'h554 == _T_12323 ? _GEN_4 : mem_1364;
  assign _GEN_9563 = 11'h555 == _T_12323 ? _GEN_4 : mem_1365;
  assign _GEN_9564 = 11'h556 == _T_12323 ? _GEN_4 : mem_1366;
  assign _GEN_9565 = 11'h557 == _T_12323 ? _GEN_4 : mem_1367;
  assign _GEN_9566 = 11'h558 == _T_12323 ? _GEN_4 : mem_1368;
  assign _GEN_9567 = 11'h559 == _T_12323 ? _GEN_4 : mem_1369;
  assign _GEN_9568 = 11'h55a == _T_12323 ? _GEN_4 : mem_1370;
  assign _GEN_9569 = 11'h55b == _T_12323 ? _GEN_4 : mem_1371;
  assign _GEN_9570 = 11'h55c == _T_12323 ? _GEN_4 : mem_1372;
  assign _GEN_9571 = 11'h55d == _T_12323 ? _GEN_4 : mem_1373;
  assign _GEN_9572 = 11'h55e == _T_12323 ? _GEN_4 : mem_1374;
  assign _GEN_9573 = 11'h55f == _T_12323 ? _GEN_4 : mem_1375;
  assign _GEN_9574 = 11'h560 == _T_12323 ? _GEN_4 : mem_1376;
  assign _GEN_9575 = 11'h561 == _T_12323 ? _GEN_4 : mem_1377;
  assign _GEN_9576 = 11'h562 == _T_12323 ? _GEN_4 : mem_1378;
  assign _GEN_9577 = 11'h563 == _T_12323 ? _GEN_4 : mem_1379;
  assign _GEN_9578 = 11'h564 == _T_12323 ? _GEN_4 : mem_1380;
  assign _GEN_9579 = 11'h565 == _T_12323 ? _GEN_4 : mem_1381;
  assign _GEN_9580 = 11'h566 == _T_12323 ? _GEN_4 : mem_1382;
  assign _GEN_9581 = 11'h567 == _T_12323 ? _GEN_4 : mem_1383;
  assign _GEN_9582 = 11'h568 == _T_12323 ? _GEN_4 : mem_1384;
  assign _GEN_9583 = 11'h569 == _T_12323 ? _GEN_4 : mem_1385;
  assign _GEN_9584 = 11'h56a == _T_12323 ? _GEN_4 : mem_1386;
  assign _GEN_9585 = 11'h56b == _T_12323 ? _GEN_4 : mem_1387;
  assign _GEN_9586 = 11'h56c == _T_12323 ? _GEN_4 : mem_1388;
  assign _GEN_9587 = 11'h56d == _T_12323 ? _GEN_4 : mem_1389;
  assign _GEN_9588 = 11'h56e == _T_12323 ? _GEN_4 : mem_1390;
  assign _GEN_9589 = 11'h56f == _T_12323 ? _GEN_4 : mem_1391;
  assign _GEN_9590 = 11'h570 == _T_12323 ? _GEN_4 : mem_1392;
  assign _GEN_9591 = 11'h571 == _T_12323 ? _GEN_4 : mem_1393;
  assign _GEN_9592 = 11'h572 == _T_12323 ? _GEN_4 : mem_1394;
  assign _GEN_9593 = 11'h573 == _T_12323 ? _GEN_4 : mem_1395;
  assign _GEN_9594 = 11'h574 == _T_12323 ? _GEN_4 : mem_1396;
  assign _GEN_9595 = 11'h575 == _T_12323 ? _GEN_4 : mem_1397;
  assign _GEN_9596 = 11'h576 == _T_12323 ? _GEN_4 : mem_1398;
  assign _GEN_9597 = 11'h577 == _T_12323 ? _GEN_4 : mem_1399;
  assign _GEN_9598 = 11'h578 == _T_12323 ? _GEN_4 : mem_1400;
  assign _GEN_9599 = 11'h579 == _T_12323 ? _GEN_4 : mem_1401;
  assign _GEN_9600 = 11'h57a == _T_12323 ? _GEN_4 : mem_1402;
  assign _GEN_9601 = 11'h57b == _T_12323 ? _GEN_4 : mem_1403;
  assign _GEN_9602 = 11'h57c == _T_12323 ? _GEN_4 : mem_1404;
  assign _GEN_9603 = 11'h57d == _T_12323 ? _GEN_4 : mem_1405;
  assign _GEN_9604 = 11'h57e == _T_12323 ? _GEN_4 : mem_1406;
  assign _GEN_9605 = 11'h57f == _T_12323 ? _GEN_4 : mem_1407;
  assign _GEN_9606 = 11'h580 == _T_12323 ? _GEN_4 : mem_1408;
  assign _GEN_9607 = 11'h581 == _T_12323 ? _GEN_4 : mem_1409;
  assign _GEN_9608 = 11'h582 == _T_12323 ? _GEN_4 : mem_1410;
  assign _GEN_9609 = 11'h583 == _T_12323 ? _GEN_4 : mem_1411;
  assign _GEN_9610 = 11'h584 == _T_12323 ? _GEN_4 : mem_1412;
  assign _GEN_9611 = 11'h585 == _T_12323 ? _GEN_4 : mem_1413;
  assign _GEN_9612 = 11'h586 == _T_12323 ? _GEN_4 : mem_1414;
  assign _GEN_9613 = 11'h587 == _T_12323 ? _GEN_4 : mem_1415;
  assign _GEN_9614 = 11'h588 == _T_12323 ? _GEN_4 : mem_1416;
  assign _GEN_9615 = 11'h589 == _T_12323 ? _GEN_4 : mem_1417;
  assign _GEN_9616 = 11'h58a == _T_12323 ? _GEN_4 : mem_1418;
  assign _GEN_9617 = 11'h58b == _T_12323 ? _GEN_4 : mem_1419;
  assign _GEN_9618 = 11'h58c == _T_12323 ? _GEN_4 : mem_1420;
  assign _GEN_9619 = 11'h58d == _T_12323 ? _GEN_4 : mem_1421;
  assign _GEN_9620 = 11'h58e == _T_12323 ? _GEN_4 : mem_1422;
  assign _GEN_9621 = 11'h58f == _T_12323 ? _GEN_4 : mem_1423;
  assign _GEN_9622 = 11'h590 == _T_12323 ? _GEN_4 : mem_1424;
  assign _GEN_9623 = 11'h591 == _T_12323 ? _GEN_4 : mem_1425;
  assign _GEN_9624 = 11'h592 == _T_12323 ? _GEN_4 : mem_1426;
  assign _GEN_9625 = 11'h593 == _T_12323 ? _GEN_4 : mem_1427;
  assign _GEN_9626 = 11'h594 == _T_12323 ? _GEN_4 : mem_1428;
  assign _GEN_9627 = 11'h595 == _T_12323 ? _GEN_4 : mem_1429;
  assign _GEN_9628 = 11'h596 == _T_12323 ? _GEN_4 : mem_1430;
  assign _GEN_9629 = 11'h597 == _T_12323 ? _GEN_4 : mem_1431;
  assign _GEN_9630 = 11'h598 == _T_12323 ? _GEN_4 : mem_1432;
  assign _GEN_9631 = 11'h599 == _T_12323 ? _GEN_4 : mem_1433;
  assign _GEN_9632 = 11'h59a == _T_12323 ? _GEN_4 : mem_1434;
  assign _GEN_9633 = 11'h59b == _T_12323 ? _GEN_4 : mem_1435;
  assign _GEN_9634 = 11'h59c == _T_12323 ? _GEN_4 : mem_1436;
  assign _GEN_9635 = 11'h59d == _T_12323 ? _GEN_4 : mem_1437;
  assign _GEN_9636 = 11'h59e == _T_12323 ? _GEN_4 : mem_1438;
  assign _GEN_9637 = 11'h59f == _T_12323 ? _GEN_4 : mem_1439;
  assign _GEN_9638 = 11'h5a0 == _T_12323 ? _GEN_4 : mem_1440;
  assign _GEN_9639 = 11'h5a1 == _T_12323 ? _GEN_4 : mem_1441;
  assign _GEN_9640 = 11'h5a2 == _T_12323 ? _GEN_4 : mem_1442;
  assign _GEN_9641 = 11'h5a3 == _T_12323 ? _GEN_4 : mem_1443;
  assign _GEN_9642 = 11'h5a4 == _T_12323 ? _GEN_4 : mem_1444;
  assign _GEN_9643 = 11'h5a5 == _T_12323 ? _GEN_4 : mem_1445;
  assign _GEN_9644 = 11'h5a6 == _T_12323 ? _GEN_4 : mem_1446;
  assign _GEN_9645 = 11'h5a7 == _T_12323 ? _GEN_4 : mem_1447;
  assign _GEN_9646 = 11'h5a8 == _T_12323 ? _GEN_4 : mem_1448;
  assign _GEN_9647 = 11'h5a9 == _T_12323 ? _GEN_4 : mem_1449;
  assign _GEN_9648 = 11'h5aa == _T_12323 ? _GEN_4 : mem_1450;
  assign _GEN_9649 = 11'h5ab == _T_12323 ? _GEN_4 : mem_1451;
  assign _GEN_9650 = 11'h5ac == _T_12323 ? _GEN_4 : mem_1452;
  assign _GEN_9651 = 11'h5ad == _T_12323 ? _GEN_4 : mem_1453;
  assign _GEN_9652 = 11'h5ae == _T_12323 ? _GEN_4 : mem_1454;
  assign _GEN_9653 = 11'h5af == _T_12323 ? _GEN_4 : mem_1455;
  assign _GEN_9654 = 11'h5b0 == _T_12323 ? _GEN_4 : mem_1456;
  assign _GEN_9655 = 11'h5b1 == _T_12323 ? _GEN_4 : mem_1457;
  assign _GEN_9656 = 11'h5b2 == _T_12323 ? _GEN_4 : mem_1458;
  assign _GEN_9657 = 11'h5b3 == _T_12323 ? _GEN_4 : mem_1459;
  assign _GEN_9658 = 11'h5b4 == _T_12323 ? _GEN_4 : mem_1460;
  assign _GEN_9659 = 11'h5b5 == _T_12323 ? _GEN_4 : mem_1461;
  assign _GEN_9660 = 11'h5b6 == _T_12323 ? _GEN_4 : mem_1462;
  assign _GEN_9661 = 11'h5b7 == _T_12323 ? _GEN_4 : mem_1463;
  assign _GEN_9662 = 11'h5b8 == _T_12323 ? _GEN_4 : mem_1464;
  assign _GEN_9663 = 11'h5b9 == _T_12323 ? _GEN_4 : mem_1465;
  assign _GEN_9664 = 11'h5ba == _T_12323 ? _GEN_4 : mem_1466;
  assign _GEN_9665 = 11'h5bb == _T_12323 ? _GEN_4 : mem_1467;
  assign _GEN_9666 = 11'h5bc == _T_12323 ? _GEN_4 : mem_1468;
  assign _GEN_9667 = 11'h5bd == _T_12323 ? _GEN_4 : mem_1469;
  assign _GEN_9668 = 11'h5be == _T_12323 ? _GEN_4 : mem_1470;
  assign _GEN_9669 = 11'h5bf == _T_12323 ? _GEN_4 : mem_1471;
  assign _GEN_9670 = 11'h5c0 == _T_12323 ? _GEN_4 : mem_1472;
  assign _GEN_9671 = 11'h5c1 == _T_12323 ? _GEN_4 : mem_1473;
  assign _GEN_9672 = 11'h5c2 == _T_12323 ? _GEN_4 : mem_1474;
  assign _GEN_9673 = 11'h5c3 == _T_12323 ? _GEN_4 : mem_1475;
  assign _GEN_9674 = 11'h5c4 == _T_12323 ? _GEN_4 : mem_1476;
  assign _GEN_9675 = 11'h5c5 == _T_12323 ? _GEN_4 : mem_1477;
  assign _GEN_9676 = 11'h5c6 == _T_12323 ? _GEN_4 : mem_1478;
  assign _GEN_9677 = 11'h5c7 == _T_12323 ? _GEN_4 : mem_1479;
  assign _GEN_9678 = 11'h5c8 == _T_12323 ? _GEN_4 : mem_1480;
  assign _GEN_9679 = 11'h5c9 == _T_12323 ? _GEN_4 : mem_1481;
  assign _GEN_9680 = 11'h5ca == _T_12323 ? _GEN_4 : mem_1482;
  assign _GEN_9681 = 11'h5cb == _T_12323 ? _GEN_4 : mem_1483;
  assign _GEN_9682 = 11'h5cc == _T_12323 ? _GEN_4 : mem_1484;
  assign _GEN_9683 = 11'h5cd == _T_12323 ? _GEN_4 : mem_1485;
  assign _GEN_9684 = 11'h5ce == _T_12323 ? _GEN_4 : mem_1486;
  assign _GEN_9685 = 11'h5cf == _T_12323 ? _GEN_4 : mem_1487;
  assign _GEN_9686 = 11'h5d0 == _T_12323 ? _GEN_4 : mem_1488;
  assign _GEN_9687 = 11'h5d1 == _T_12323 ? _GEN_4 : mem_1489;
  assign _GEN_9688 = 11'h5d2 == _T_12323 ? _GEN_4 : mem_1490;
  assign _GEN_9689 = 11'h5d3 == _T_12323 ? _GEN_4 : mem_1491;
  assign _GEN_9690 = 11'h5d4 == _T_12323 ? _GEN_4 : mem_1492;
  assign _GEN_9691 = 11'h5d5 == _T_12323 ? _GEN_4 : mem_1493;
  assign _GEN_9692 = 11'h5d6 == _T_12323 ? _GEN_4 : mem_1494;
  assign _GEN_9693 = 11'h5d7 == _T_12323 ? _GEN_4 : mem_1495;
  assign _GEN_9694 = 11'h5d8 == _T_12323 ? _GEN_4 : mem_1496;
  assign _GEN_9695 = 11'h5d9 == _T_12323 ? _GEN_4 : mem_1497;
  assign _GEN_9696 = 11'h5da == _T_12323 ? _GEN_4 : mem_1498;
  assign _GEN_9697 = 11'h5db == _T_12323 ? _GEN_4 : mem_1499;
  assign _GEN_9698 = 11'h5dc == _T_12323 ? _GEN_4 : mem_1500;
  assign _GEN_9699 = 11'h5dd == _T_12323 ? _GEN_4 : mem_1501;
  assign _GEN_9700 = 11'h5de == _T_12323 ? _GEN_4 : mem_1502;
  assign _GEN_9701 = 11'h5df == _T_12323 ? _GEN_4 : mem_1503;
  assign _GEN_9702 = 11'h5e0 == _T_12323 ? _GEN_4 : mem_1504;
  assign _GEN_9703 = 11'h5e1 == _T_12323 ? _GEN_4 : mem_1505;
  assign _GEN_9704 = 11'h5e2 == _T_12323 ? _GEN_4 : mem_1506;
  assign _GEN_9705 = 11'h5e3 == _T_12323 ? _GEN_4 : mem_1507;
  assign _GEN_9706 = 11'h5e4 == _T_12323 ? _GEN_4 : mem_1508;
  assign _GEN_9707 = 11'h5e5 == _T_12323 ? _GEN_4 : mem_1509;
  assign _GEN_9708 = 11'h5e6 == _T_12323 ? _GEN_4 : mem_1510;
  assign _GEN_9709 = 11'h5e7 == _T_12323 ? _GEN_4 : mem_1511;
  assign _GEN_9710 = 11'h5e8 == _T_12323 ? _GEN_4 : mem_1512;
  assign _GEN_9711 = 11'h5e9 == _T_12323 ? _GEN_4 : mem_1513;
  assign _GEN_9712 = 11'h5ea == _T_12323 ? _GEN_4 : mem_1514;
  assign _GEN_9713 = 11'h5eb == _T_12323 ? _GEN_4 : mem_1515;
  assign _GEN_9714 = 11'h5ec == _T_12323 ? _GEN_4 : mem_1516;
  assign _GEN_9715 = 11'h5ed == _T_12323 ? _GEN_4 : mem_1517;
  assign _GEN_9716 = 11'h5ee == _T_12323 ? _GEN_4 : mem_1518;
  assign _GEN_9717 = 11'h5ef == _T_12323 ? _GEN_4 : mem_1519;
  assign _GEN_9718 = 11'h5f0 == _T_12323 ? _GEN_4 : mem_1520;
  assign _GEN_9719 = 11'h5f1 == _T_12323 ? _GEN_4 : mem_1521;
  assign _GEN_9720 = 11'h5f2 == _T_12323 ? _GEN_4 : mem_1522;
  assign _GEN_9721 = 11'h5f3 == _T_12323 ? _GEN_4 : mem_1523;
  assign _GEN_9722 = 11'h5f4 == _T_12323 ? _GEN_4 : mem_1524;
  assign _GEN_9723 = 11'h5f5 == _T_12323 ? _GEN_4 : mem_1525;
  assign _GEN_9724 = 11'h5f6 == _T_12323 ? _GEN_4 : mem_1526;
  assign _GEN_9725 = 11'h5f7 == _T_12323 ? _GEN_4 : mem_1527;
  assign _GEN_9726 = 11'h5f8 == _T_12323 ? _GEN_4 : mem_1528;
  assign _GEN_9727 = 11'h5f9 == _T_12323 ? _GEN_4 : mem_1529;
  assign _GEN_9728 = 11'h5fa == _T_12323 ? _GEN_4 : mem_1530;
  assign _GEN_9729 = 11'h5fb == _T_12323 ? _GEN_4 : mem_1531;
  assign _GEN_9730 = 11'h5fc == _T_12323 ? _GEN_4 : mem_1532;
  assign _GEN_9731 = 11'h5fd == _T_12323 ? _GEN_4 : mem_1533;
  assign _GEN_9732 = 11'h5fe == _T_12323 ? _GEN_4 : mem_1534;
  assign _GEN_9733 = 11'h5ff == _T_12323 ? _GEN_4 : mem_1535;
  assign _GEN_9734 = 11'h600 == _T_12323 ? _GEN_4 : mem_1536;
  assign _GEN_9735 = 11'h601 == _T_12323 ? _GEN_4 : mem_1537;
  assign _GEN_9736 = 11'h602 == _T_12323 ? _GEN_4 : mem_1538;
  assign _GEN_9737 = 11'h603 == _T_12323 ? _GEN_4 : mem_1539;
  assign _GEN_9738 = 11'h604 == _T_12323 ? _GEN_4 : mem_1540;
  assign _GEN_9739 = 11'h605 == _T_12323 ? _GEN_4 : mem_1541;
  assign _GEN_9740 = 11'h606 == _T_12323 ? _GEN_4 : mem_1542;
  assign _GEN_9741 = 11'h607 == _T_12323 ? _GEN_4 : mem_1543;
  assign _GEN_9742 = 11'h608 == _T_12323 ? _GEN_4 : mem_1544;
  assign _GEN_9743 = 11'h609 == _T_12323 ? _GEN_4 : mem_1545;
  assign _GEN_9744 = 11'h60a == _T_12323 ? _GEN_4 : mem_1546;
  assign _GEN_9745 = 11'h60b == _T_12323 ? _GEN_4 : mem_1547;
  assign _GEN_9746 = 11'h60c == _T_12323 ? _GEN_4 : mem_1548;
  assign _GEN_9747 = 11'h60d == _T_12323 ? _GEN_4 : mem_1549;
  assign _GEN_9748 = 11'h60e == _T_12323 ? _GEN_4 : mem_1550;
  assign _GEN_9749 = 11'h60f == _T_12323 ? _GEN_4 : mem_1551;
  assign _GEN_9750 = 11'h610 == _T_12323 ? _GEN_4 : mem_1552;
  assign _GEN_9751 = 11'h611 == _T_12323 ? _GEN_4 : mem_1553;
  assign _GEN_9752 = 11'h612 == _T_12323 ? _GEN_4 : mem_1554;
  assign _GEN_9753 = 11'h613 == _T_12323 ? _GEN_4 : mem_1555;
  assign _GEN_9754 = 11'h614 == _T_12323 ? _GEN_4 : mem_1556;
  assign _GEN_9755 = 11'h615 == _T_12323 ? _GEN_4 : mem_1557;
  assign _GEN_9756 = 11'h616 == _T_12323 ? _GEN_4 : mem_1558;
  assign _GEN_9757 = 11'h617 == _T_12323 ? _GEN_4 : mem_1559;
  assign _GEN_9758 = 11'h618 == _T_12323 ? _GEN_4 : mem_1560;
  assign _GEN_9759 = 11'h619 == _T_12323 ? _GEN_4 : mem_1561;
  assign _GEN_9760 = 11'h61a == _T_12323 ? _GEN_4 : mem_1562;
  assign _GEN_9761 = 11'h61b == _T_12323 ? _GEN_4 : mem_1563;
  assign _GEN_9762 = 11'h61c == _T_12323 ? _GEN_4 : mem_1564;
  assign _GEN_9763 = 11'h61d == _T_12323 ? _GEN_4 : mem_1565;
  assign _GEN_9764 = 11'h61e == _T_12323 ? _GEN_4 : mem_1566;
  assign _GEN_9765 = 11'h61f == _T_12323 ? _GEN_4 : mem_1567;
  assign _GEN_9766 = 11'h620 == _T_12323 ? _GEN_4 : mem_1568;
  assign _GEN_9767 = 11'h621 == _T_12323 ? _GEN_4 : mem_1569;
  assign _GEN_9768 = 11'h622 == _T_12323 ? _GEN_4 : mem_1570;
  assign _GEN_9769 = 11'h623 == _T_12323 ? _GEN_4 : mem_1571;
  assign _GEN_9770 = 11'h624 == _T_12323 ? _GEN_4 : mem_1572;
  assign _GEN_9771 = 11'h625 == _T_12323 ? _GEN_4 : mem_1573;
  assign _GEN_9772 = 11'h626 == _T_12323 ? _GEN_4 : mem_1574;
  assign _GEN_9773 = 11'h627 == _T_12323 ? _GEN_4 : mem_1575;
  assign _GEN_9774 = 11'h628 == _T_12323 ? _GEN_4 : mem_1576;
  assign _GEN_9775 = 11'h629 == _T_12323 ? _GEN_4 : mem_1577;
  assign _GEN_9776 = 11'h62a == _T_12323 ? _GEN_4 : mem_1578;
  assign _GEN_9777 = 11'h62b == _T_12323 ? _GEN_4 : mem_1579;
  assign _GEN_9778 = 11'h62c == _T_12323 ? _GEN_4 : mem_1580;
  assign _GEN_9779 = 11'h62d == _T_12323 ? _GEN_4 : mem_1581;
  assign _GEN_9780 = 11'h62e == _T_12323 ? _GEN_4 : mem_1582;
  assign _GEN_9781 = 11'h62f == _T_12323 ? _GEN_4 : mem_1583;
  assign _GEN_9782 = 11'h630 == _T_12323 ? _GEN_4 : mem_1584;
  assign _GEN_9783 = 11'h631 == _T_12323 ? _GEN_4 : mem_1585;
  assign _GEN_9784 = 11'h632 == _T_12323 ? _GEN_4 : mem_1586;
  assign _GEN_9785 = 11'h633 == _T_12323 ? _GEN_4 : mem_1587;
  assign _GEN_9786 = 11'h634 == _T_12323 ? _GEN_4 : mem_1588;
  assign _GEN_9787 = 11'h635 == _T_12323 ? _GEN_4 : mem_1589;
  assign _GEN_9788 = 11'h636 == _T_12323 ? _GEN_4 : mem_1590;
  assign _GEN_9789 = 11'h637 == _T_12323 ? _GEN_4 : mem_1591;
  assign _GEN_9790 = 11'h638 == _T_12323 ? _GEN_4 : mem_1592;
  assign _GEN_9791 = 11'h639 == _T_12323 ? _GEN_4 : mem_1593;
  assign _GEN_9792 = 11'h63a == _T_12323 ? _GEN_4 : mem_1594;
  assign _GEN_9793 = 11'h63b == _T_12323 ? _GEN_4 : mem_1595;
  assign _GEN_9794 = 11'h63c == _T_12323 ? _GEN_4 : mem_1596;
  assign _GEN_9795 = 11'h63d == _T_12323 ? _GEN_4 : mem_1597;
  assign _GEN_9796 = 11'h63e == _T_12323 ? _GEN_4 : mem_1598;
  assign _GEN_9797 = 11'h63f == _T_12323 ? _GEN_4 : mem_1599;
  assign _GEN_9798 = 11'h640 == _T_12323 ? _GEN_4 : mem_1600;
  assign _GEN_9799 = 11'h641 == _T_12323 ? _GEN_4 : mem_1601;
  assign _GEN_9800 = 11'h642 == _T_12323 ? _GEN_4 : mem_1602;
  assign _GEN_9801 = 11'h643 == _T_12323 ? _GEN_4 : mem_1603;
  assign _GEN_9802 = 11'h644 == _T_12323 ? _GEN_4 : mem_1604;
  assign _GEN_9803 = 11'h645 == _T_12323 ? _GEN_4 : mem_1605;
  assign _GEN_9804 = 11'h646 == _T_12323 ? _GEN_4 : mem_1606;
  assign _GEN_9805 = 11'h647 == _T_12323 ? _GEN_4 : mem_1607;
  assign _GEN_9806 = 11'h648 == _T_12323 ? _GEN_4 : mem_1608;
  assign _GEN_9807 = 11'h649 == _T_12323 ? _GEN_4 : mem_1609;
  assign _GEN_9808 = 11'h64a == _T_12323 ? _GEN_4 : mem_1610;
  assign _GEN_9809 = 11'h64b == _T_12323 ? _GEN_4 : mem_1611;
  assign _GEN_9810 = 11'h64c == _T_12323 ? _GEN_4 : mem_1612;
  assign _GEN_9811 = 11'h64d == _T_12323 ? _GEN_4 : mem_1613;
  assign _GEN_9812 = 11'h64e == _T_12323 ? _GEN_4 : mem_1614;
  assign _GEN_9813 = 11'h64f == _T_12323 ? _GEN_4 : mem_1615;
  assign _GEN_9814 = 11'h650 == _T_12323 ? _GEN_4 : mem_1616;
  assign _GEN_9815 = 11'h651 == _T_12323 ? _GEN_4 : mem_1617;
  assign _GEN_9816 = 11'h652 == _T_12323 ? _GEN_4 : mem_1618;
  assign _GEN_9817 = 11'h653 == _T_12323 ? _GEN_4 : mem_1619;
  assign _GEN_9818 = 11'h654 == _T_12323 ? _GEN_4 : mem_1620;
  assign _GEN_9819 = 11'h655 == _T_12323 ? _GEN_4 : mem_1621;
  assign _GEN_9820 = 11'h656 == _T_12323 ? _GEN_4 : mem_1622;
  assign _GEN_9821 = 11'h657 == _T_12323 ? _GEN_4 : mem_1623;
  assign _GEN_9822 = 11'h658 == _T_12323 ? _GEN_4 : mem_1624;
  assign _GEN_9823 = 11'h659 == _T_12323 ? _GEN_4 : mem_1625;
  assign _GEN_9824 = 11'h65a == _T_12323 ? _GEN_4 : mem_1626;
  assign _GEN_9825 = 11'h65b == _T_12323 ? _GEN_4 : mem_1627;
  assign _GEN_9826 = 11'h65c == _T_12323 ? _GEN_4 : mem_1628;
  assign _GEN_9827 = 11'h65d == _T_12323 ? _GEN_4 : mem_1629;
  assign _GEN_9828 = 11'h65e == _T_12323 ? _GEN_4 : mem_1630;
  assign _GEN_9829 = 11'h65f == _T_12323 ? _GEN_4 : mem_1631;
  assign _GEN_9830 = 11'h660 == _T_12323 ? _GEN_4 : mem_1632;
  assign _GEN_9831 = 11'h661 == _T_12323 ? _GEN_4 : mem_1633;
  assign _GEN_9832 = 11'h662 == _T_12323 ? _GEN_4 : mem_1634;
  assign _GEN_9833 = 11'h663 == _T_12323 ? _GEN_4 : mem_1635;
  assign _GEN_9834 = 11'h664 == _T_12323 ? _GEN_4 : mem_1636;
  assign _GEN_9835 = 11'h665 == _T_12323 ? _GEN_4 : mem_1637;
  assign _GEN_9836 = 11'h666 == _T_12323 ? _GEN_4 : mem_1638;
  assign _GEN_9837 = 11'h667 == _T_12323 ? _GEN_4 : mem_1639;
  assign _GEN_9838 = 11'h668 == _T_12323 ? _GEN_4 : mem_1640;
  assign _GEN_9839 = 11'h669 == _T_12323 ? _GEN_4 : mem_1641;
  assign _GEN_9840 = 11'h66a == _T_12323 ? _GEN_4 : mem_1642;
  assign _GEN_9841 = 11'h66b == _T_12323 ? _GEN_4 : mem_1643;
  assign _GEN_9842 = 11'h66c == _T_12323 ? _GEN_4 : mem_1644;
  assign _GEN_9843 = 11'h66d == _T_12323 ? _GEN_4 : mem_1645;
  assign _GEN_9844 = 11'h66e == _T_12323 ? _GEN_4 : mem_1646;
  assign _GEN_9845 = 11'h66f == _T_12323 ? _GEN_4 : mem_1647;
  assign _GEN_9846 = 11'h670 == _T_12323 ? _GEN_4 : mem_1648;
  assign _GEN_9847 = 11'h671 == _T_12323 ? _GEN_4 : mem_1649;
  assign _GEN_9848 = 11'h672 == _T_12323 ? _GEN_4 : mem_1650;
  assign _GEN_9849 = 11'h673 == _T_12323 ? _GEN_4 : mem_1651;
  assign _GEN_9850 = 11'h674 == _T_12323 ? _GEN_4 : mem_1652;
  assign _GEN_9851 = 11'h675 == _T_12323 ? _GEN_4 : mem_1653;
  assign _GEN_9852 = 11'h676 == _T_12323 ? _GEN_4 : mem_1654;
  assign _GEN_9853 = 11'h677 == _T_12323 ? _GEN_4 : mem_1655;
  assign _GEN_9854 = 11'h678 == _T_12323 ? _GEN_4 : mem_1656;
  assign _GEN_9855 = 11'h679 == _T_12323 ? _GEN_4 : mem_1657;
  assign _GEN_9856 = 11'h67a == _T_12323 ? _GEN_4 : mem_1658;
  assign _GEN_9857 = 11'h67b == _T_12323 ? _GEN_4 : mem_1659;
  assign _GEN_9858 = 11'h67c == _T_12323 ? _GEN_4 : mem_1660;
  assign _GEN_9859 = 11'h67d == _T_12323 ? _GEN_4 : mem_1661;
  assign _GEN_9860 = 11'h67e == _T_12323 ? _GEN_4 : mem_1662;
  assign _GEN_9861 = 11'h67f == _T_12323 ? _GEN_4 : mem_1663;
  assign _GEN_9862 = 11'h680 == _T_12323 ? _GEN_4 : mem_1664;
  assign _GEN_9863 = 11'h681 == _T_12323 ? _GEN_4 : mem_1665;
  assign _GEN_9864 = 11'h682 == _T_12323 ? _GEN_4 : mem_1666;
  assign _GEN_9865 = 11'h683 == _T_12323 ? _GEN_4 : mem_1667;
  assign _GEN_9866 = 11'h684 == _T_12323 ? _GEN_4 : mem_1668;
  assign _GEN_9867 = 11'h685 == _T_12323 ? _GEN_4 : mem_1669;
  assign _GEN_9868 = 11'h686 == _T_12323 ? _GEN_4 : mem_1670;
  assign _GEN_9869 = 11'h687 == _T_12323 ? _GEN_4 : mem_1671;
  assign _GEN_9870 = 11'h688 == _T_12323 ? _GEN_4 : mem_1672;
  assign _GEN_9871 = 11'h689 == _T_12323 ? _GEN_4 : mem_1673;
  assign _GEN_9872 = 11'h68a == _T_12323 ? _GEN_4 : mem_1674;
  assign _GEN_9873 = 11'h68b == _T_12323 ? _GEN_4 : mem_1675;
  assign _GEN_9874 = 11'h68c == _T_12323 ? _GEN_4 : mem_1676;
  assign _GEN_9875 = 11'h68d == _T_12323 ? _GEN_4 : mem_1677;
  assign _GEN_9876 = 11'h68e == _T_12323 ? _GEN_4 : mem_1678;
  assign _GEN_9877 = 11'h68f == _T_12323 ? _GEN_4 : mem_1679;
  assign _GEN_9878 = 11'h690 == _T_12323 ? _GEN_4 : mem_1680;
  assign _GEN_9879 = 11'h691 == _T_12323 ? _GEN_4 : mem_1681;
  assign _GEN_9880 = 11'h692 == _T_12323 ? _GEN_4 : mem_1682;
  assign _GEN_9881 = 11'h693 == _T_12323 ? _GEN_4 : mem_1683;
  assign _GEN_9882 = 11'h694 == _T_12323 ? _GEN_4 : mem_1684;
  assign _GEN_9883 = 11'h695 == _T_12323 ? _GEN_4 : mem_1685;
  assign _GEN_9884 = 11'h696 == _T_12323 ? _GEN_4 : mem_1686;
  assign _GEN_9885 = 11'h697 == _T_12323 ? _GEN_4 : mem_1687;
  assign _GEN_9886 = 11'h698 == _T_12323 ? _GEN_4 : mem_1688;
  assign _GEN_9887 = 11'h699 == _T_12323 ? _GEN_4 : mem_1689;
  assign _GEN_9888 = 11'h69a == _T_12323 ? _GEN_4 : mem_1690;
  assign _GEN_9889 = 11'h69b == _T_12323 ? _GEN_4 : mem_1691;
  assign _GEN_9890 = 11'h69c == _T_12323 ? _GEN_4 : mem_1692;
  assign _GEN_9891 = 11'h69d == _T_12323 ? _GEN_4 : mem_1693;
  assign _GEN_9892 = 11'h69e == _T_12323 ? _GEN_4 : mem_1694;
  assign _GEN_9893 = 11'h69f == _T_12323 ? _GEN_4 : mem_1695;
  assign _GEN_9894 = 11'h6a0 == _T_12323 ? _GEN_4 : mem_1696;
  assign _GEN_9895 = 11'h6a1 == _T_12323 ? _GEN_4 : mem_1697;
  assign _GEN_9896 = 11'h6a2 == _T_12323 ? _GEN_4 : mem_1698;
  assign _GEN_9897 = 11'h6a3 == _T_12323 ? _GEN_4 : mem_1699;
  assign _GEN_9898 = 11'h6a4 == _T_12323 ? _GEN_4 : mem_1700;
  assign _GEN_9899 = 11'h6a5 == _T_12323 ? _GEN_4 : mem_1701;
  assign _GEN_9900 = 11'h6a6 == _T_12323 ? _GEN_4 : mem_1702;
  assign _GEN_9901 = 11'h6a7 == _T_12323 ? _GEN_4 : mem_1703;
  assign _GEN_9902 = 11'h6a8 == _T_12323 ? _GEN_4 : mem_1704;
  assign _GEN_9903 = 11'h6a9 == _T_12323 ? _GEN_4 : mem_1705;
  assign _GEN_9904 = 11'h6aa == _T_12323 ? _GEN_4 : mem_1706;
  assign _GEN_9905 = 11'h6ab == _T_12323 ? _GEN_4 : mem_1707;
  assign _GEN_9906 = 11'h6ac == _T_12323 ? _GEN_4 : mem_1708;
  assign _GEN_9907 = 11'h6ad == _T_12323 ? _GEN_4 : mem_1709;
  assign _GEN_9908 = 11'h6ae == _T_12323 ? _GEN_4 : mem_1710;
  assign _GEN_9909 = 11'h6af == _T_12323 ? _GEN_4 : mem_1711;
  assign _GEN_9910 = 11'h6b0 == _T_12323 ? _GEN_4 : mem_1712;
  assign _GEN_9911 = 11'h6b1 == _T_12323 ? _GEN_4 : mem_1713;
  assign _GEN_9912 = 11'h6b2 == _T_12323 ? _GEN_4 : mem_1714;
  assign _GEN_9913 = 11'h6b3 == _T_12323 ? _GEN_4 : mem_1715;
  assign _GEN_9914 = 11'h6b4 == _T_12323 ? _GEN_4 : mem_1716;
  assign _GEN_9915 = 11'h6b5 == _T_12323 ? _GEN_4 : mem_1717;
  assign _GEN_9916 = 11'h6b6 == _T_12323 ? _GEN_4 : mem_1718;
  assign _GEN_9917 = 11'h6b7 == _T_12323 ? _GEN_4 : mem_1719;
  assign _GEN_9918 = 11'h6b8 == _T_12323 ? _GEN_4 : mem_1720;
  assign _GEN_9919 = 11'h6b9 == _T_12323 ? _GEN_4 : mem_1721;
  assign _GEN_9920 = 11'h6ba == _T_12323 ? _GEN_4 : mem_1722;
  assign _GEN_9921 = 11'h6bb == _T_12323 ? _GEN_4 : mem_1723;
  assign _GEN_9922 = 11'h6bc == _T_12323 ? _GEN_4 : mem_1724;
  assign _GEN_9923 = 11'h6bd == _T_12323 ? _GEN_4 : mem_1725;
  assign _GEN_9924 = 11'h6be == _T_12323 ? _GEN_4 : mem_1726;
  assign _GEN_9925 = 11'h6bf == _T_12323 ? _GEN_4 : mem_1727;
  assign _GEN_9926 = 11'h6c0 == _T_12323 ? _GEN_4 : mem_1728;
  assign _GEN_9927 = 11'h6c1 == _T_12323 ? _GEN_4 : mem_1729;
  assign _GEN_9928 = 11'h6c2 == _T_12323 ? _GEN_4 : mem_1730;
  assign _GEN_9929 = 11'h6c3 == _T_12323 ? _GEN_4 : mem_1731;
  assign _GEN_9930 = 11'h6c4 == _T_12323 ? _GEN_4 : mem_1732;
  assign _GEN_9931 = 11'h6c5 == _T_12323 ? _GEN_4 : mem_1733;
  assign _GEN_9932 = 11'h6c6 == _T_12323 ? _GEN_4 : mem_1734;
  assign _GEN_9933 = 11'h6c7 == _T_12323 ? _GEN_4 : mem_1735;
  assign _GEN_9934 = 11'h6c8 == _T_12323 ? _GEN_4 : mem_1736;
  assign _GEN_9935 = 11'h6c9 == _T_12323 ? _GEN_4 : mem_1737;
  assign _GEN_9936 = 11'h6ca == _T_12323 ? _GEN_4 : mem_1738;
  assign _GEN_9937 = 11'h6cb == _T_12323 ? _GEN_4 : mem_1739;
  assign _GEN_9938 = 11'h6cc == _T_12323 ? _GEN_4 : mem_1740;
  assign _GEN_9939 = 11'h6cd == _T_12323 ? _GEN_4 : mem_1741;
  assign _GEN_9940 = 11'h6ce == _T_12323 ? _GEN_4 : mem_1742;
  assign _GEN_9941 = 11'h6cf == _T_12323 ? _GEN_4 : mem_1743;
  assign _GEN_9942 = 11'h6d0 == _T_12323 ? _GEN_4 : mem_1744;
  assign _GEN_9943 = 11'h6d1 == _T_12323 ? _GEN_4 : mem_1745;
  assign _GEN_9944 = 11'h6d2 == _T_12323 ? _GEN_4 : mem_1746;
  assign _GEN_9945 = 11'h6d3 == _T_12323 ? _GEN_4 : mem_1747;
  assign _GEN_9946 = 11'h6d4 == _T_12323 ? _GEN_4 : mem_1748;
  assign _GEN_9947 = 11'h6d5 == _T_12323 ? _GEN_4 : mem_1749;
  assign _GEN_9948 = 11'h6d6 == _T_12323 ? _GEN_4 : mem_1750;
  assign _GEN_9949 = 11'h6d7 == _T_12323 ? _GEN_4 : mem_1751;
  assign _GEN_9950 = 11'h6d8 == _T_12323 ? _GEN_4 : mem_1752;
  assign _GEN_9951 = 11'h6d9 == _T_12323 ? _GEN_4 : mem_1753;
  assign _GEN_9952 = 11'h6da == _T_12323 ? _GEN_4 : mem_1754;
  assign _GEN_9953 = 11'h6db == _T_12323 ? _GEN_4 : mem_1755;
  assign _GEN_9954 = 11'h6dc == _T_12323 ? _GEN_4 : mem_1756;
  assign _GEN_9955 = 11'h6dd == _T_12323 ? _GEN_4 : mem_1757;
  assign _GEN_9956 = 11'h6de == _T_12323 ? _GEN_4 : mem_1758;
  assign _GEN_9957 = 11'h6df == _T_12323 ? _GEN_4 : mem_1759;
  assign _GEN_9958 = 11'h6e0 == _T_12323 ? _GEN_4 : mem_1760;
  assign _GEN_9959 = 11'h6e1 == _T_12323 ? _GEN_4 : mem_1761;
  assign _GEN_9960 = 11'h6e2 == _T_12323 ? _GEN_4 : mem_1762;
  assign _GEN_9961 = 11'h6e3 == _T_12323 ? _GEN_4 : mem_1763;
  assign _GEN_9962 = 11'h6e4 == _T_12323 ? _GEN_4 : mem_1764;
  assign _GEN_9963 = 11'h6e5 == _T_12323 ? _GEN_4 : mem_1765;
  assign _GEN_9964 = 11'h6e6 == _T_12323 ? _GEN_4 : mem_1766;
  assign _GEN_9965 = 11'h6e7 == _T_12323 ? _GEN_4 : mem_1767;
  assign _GEN_9966 = 11'h6e8 == _T_12323 ? _GEN_4 : mem_1768;
  assign _GEN_9967 = 11'h6e9 == _T_12323 ? _GEN_4 : mem_1769;
  assign _GEN_9968 = 11'h6ea == _T_12323 ? _GEN_4 : mem_1770;
  assign _GEN_9969 = 11'h6eb == _T_12323 ? _GEN_4 : mem_1771;
  assign _GEN_9970 = 11'h6ec == _T_12323 ? _GEN_4 : mem_1772;
  assign _GEN_9971 = 11'h6ed == _T_12323 ? _GEN_4 : mem_1773;
  assign _GEN_9972 = 11'h6ee == _T_12323 ? _GEN_4 : mem_1774;
  assign _GEN_9973 = 11'h6ef == _T_12323 ? _GEN_4 : mem_1775;
  assign _GEN_9974 = 11'h6f0 == _T_12323 ? _GEN_4 : mem_1776;
  assign _GEN_9975 = 11'h6f1 == _T_12323 ? _GEN_4 : mem_1777;
  assign _GEN_9976 = 11'h6f2 == _T_12323 ? _GEN_4 : mem_1778;
  assign _GEN_9977 = 11'h6f3 == _T_12323 ? _GEN_4 : mem_1779;
  assign _GEN_9978 = 11'h6f4 == _T_12323 ? _GEN_4 : mem_1780;
  assign _GEN_9979 = 11'h6f5 == _T_12323 ? _GEN_4 : mem_1781;
  assign _GEN_9980 = 11'h6f6 == _T_12323 ? _GEN_4 : mem_1782;
  assign _GEN_9981 = 11'h6f7 == _T_12323 ? _GEN_4 : mem_1783;
  assign _GEN_9982 = 11'h6f8 == _T_12323 ? _GEN_4 : mem_1784;
  assign _GEN_9983 = 11'h6f9 == _T_12323 ? _GEN_4 : mem_1785;
  assign _GEN_9984 = 11'h6fa == _T_12323 ? _GEN_4 : mem_1786;
  assign _GEN_9985 = 11'h6fb == _T_12323 ? _GEN_4 : mem_1787;
  assign _GEN_9986 = 11'h6fc == _T_12323 ? _GEN_4 : mem_1788;
  assign _GEN_9987 = 11'h6fd == _T_12323 ? _GEN_4 : mem_1789;
  assign _GEN_9988 = 11'h6fe == _T_12323 ? _GEN_4 : mem_1790;
  assign _GEN_9989 = 11'h6ff == _T_12323 ? _GEN_4 : mem_1791;
  assign _GEN_9990 = 11'h700 == _T_12323 ? _GEN_4 : mem_1792;
  assign _GEN_9991 = 11'h701 == _T_12323 ? _GEN_4 : mem_1793;
  assign _GEN_9992 = 11'h702 == _T_12323 ? _GEN_4 : mem_1794;
  assign _GEN_9993 = 11'h703 == _T_12323 ? _GEN_4 : mem_1795;
  assign _GEN_9994 = 11'h704 == _T_12323 ? _GEN_4 : mem_1796;
  assign _GEN_9995 = 11'h705 == _T_12323 ? _GEN_4 : mem_1797;
  assign _GEN_9996 = 11'h706 == _T_12323 ? _GEN_4 : mem_1798;
  assign _GEN_9997 = 11'h707 == _T_12323 ? _GEN_4 : mem_1799;
  assign _GEN_9998 = 11'h708 == _T_12323 ? _GEN_4 : mem_1800;
  assign _GEN_9999 = 11'h709 == _T_12323 ? _GEN_4 : mem_1801;
  assign _GEN_10000 = 11'h70a == _T_12323 ? _GEN_4 : mem_1802;
  assign _GEN_10001 = 11'h70b == _T_12323 ? _GEN_4 : mem_1803;
  assign _GEN_10002 = 11'h70c == _T_12323 ? _GEN_4 : mem_1804;
  assign _GEN_10003 = 11'h70d == _T_12323 ? _GEN_4 : mem_1805;
  assign _GEN_10004 = 11'h70e == _T_12323 ? _GEN_4 : mem_1806;
  assign _GEN_10005 = 11'h70f == _T_12323 ? _GEN_4 : mem_1807;
  assign _GEN_10006 = 11'h710 == _T_12323 ? _GEN_4 : mem_1808;
  assign _GEN_10007 = 11'h711 == _T_12323 ? _GEN_4 : mem_1809;
  assign _GEN_10008 = 11'h712 == _T_12323 ? _GEN_4 : mem_1810;
  assign _GEN_10009 = 11'h713 == _T_12323 ? _GEN_4 : mem_1811;
  assign _GEN_10010 = 11'h714 == _T_12323 ? _GEN_4 : mem_1812;
  assign _GEN_10011 = 11'h715 == _T_12323 ? _GEN_4 : mem_1813;
  assign _GEN_10012 = 11'h716 == _T_12323 ? _GEN_4 : mem_1814;
  assign _GEN_10013 = 11'h717 == _T_12323 ? _GEN_4 : mem_1815;
  assign _GEN_10014 = 11'h718 == _T_12323 ? _GEN_4 : mem_1816;
  assign _GEN_10015 = 11'h719 == _T_12323 ? _GEN_4 : mem_1817;
  assign _GEN_10016 = 11'h71a == _T_12323 ? _GEN_4 : mem_1818;
  assign _GEN_10017 = 11'h71b == _T_12323 ? _GEN_4 : mem_1819;
  assign _GEN_10018 = 11'h71c == _T_12323 ? _GEN_4 : mem_1820;
  assign _GEN_10019 = 11'h71d == _T_12323 ? _GEN_4 : mem_1821;
  assign _GEN_10020 = 11'h71e == _T_12323 ? _GEN_4 : mem_1822;
  assign _GEN_10021 = 11'h71f == _T_12323 ? _GEN_4 : mem_1823;
  assign _GEN_10022 = 11'h720 == _T_12323 ? _GEN_4 : mem_1824;
  assign _GEN_10023 = 11'h721 == _T_12323 ? _GEN_4 : mem_1825;
  assign _GEN_10024 = 11'h722 == _T_12323 ? _GEN_4 : mem_1826;
  assign _GEN_10025 = 11'h723 == _T_12323 ? _GEN_4 : mem_1827;
  assign _GEN_10026 = 11'h724 == _T_12323 ? _GEN_4 : mem_1828;
  assign _GEN_10027 = 11'h725 == _T_12323 ? _GEN_4 : mem_1829;
  assign _GEN_10028 = 11'h726 == _T_12323 ? _GEN_4 : mem_1830;
  assign _GEN_10029 = 11'h727 == _T_12323 ? _GEN_4 : mem_1831;
  assign _GEN_10030 = 11'h728 == _T_12323 ? _GEN_4 : mem_1832;
  assign _GEN_10031 = 11'h729 == _T_12323 ? _GEN_4 : mem_1833;
  assign _GEN_10032 = 11'h72a == _T_12323 ? _GEN_4 : mem_1834;
  assign _GEN_10033 = 11'h72b == _T_12323 ? _GEN_4 : mem_1835;
  assign _GEN_10034 = 11'h72c == _T_12323 ? _GEN_4 : mem_1836;
  assign _GEN_10035 = 11'h72d == _T_12323 ? _GEN_4 : mem_1837;
  assign _GEN_10036 = 11'h72e == _T_12323 ? _GEN_4 : mem_1838;
  assign _GEN_10037 = 11'h72f == _T_12323 ? _GEN_4 : mem_1839;
  assign _GEN_10038 = 11'h730 == _T_12323 ? _GEN_4 : mem_1840;
  assign _GEN_10039 = 11'h731 == _T_12323 ? _GEN_4 : mem_1841;
  assign _GEN_10040 = 11'h732 == _T_12323 ? _GEN_4 : mem_1842;
  assign _GEN_10041 = 11'h733 == _T_12323 ? _GEN_4 : mem_1843;
  assign _GEN_10042 = 11'h734 == _T_12323 ? _GEN_4 : mem_1844;
  assign _GEN_10043 = 11'h735 == _T_12323 ? _GEN_4 : mem_1845;
  assign _GEN_10044 = 11'h736 == _T_12323 ? _GEN_4 : mem_1846;
  assign _GEN_10045 = 11'h737 == _T_12323 ? _GEN_4 : mem_1847;
  assign _GEN_10046 = 11'h738 == _T_12323 ? _GEN_4 : mem_1848;
  assign _GEN_10047 = 11'h739 == _T_12323 ? _GEN_4 : mem_1849;
  assign _GEN_10048 = 11'h73a == _T_12323 ? _GEN_4 : mem_1850;
  assign _GEN_10049 = 11'h73b == _T_12323 ? _GEN_4 : mem_1851;
  assign _GEN_10050 = 11'h73c == _T_12323 ? _GEN_4 : mem_1852;
  assign _GEN_10051 = 11'h73d == _T_12323 ? _GEN_4 : mem_1853;
  assign _GEN_10052 = 11'h73e == _T_12323 ? _GEN_4 : mem_1854;
  assign _GEN_10053 = 11'h73f == _T_12323 ? _GEN_4 : mem_1855;
  assign _GEN_10054 = 11'h740 == _T_12323 ? _GEN_4 : mem_1856;
  assign _GEN_10055 = 11'h741 == _T_12323 ? _GEN_4 : mem_1857;
  assign _GEN_10056 = 11'h742 == _T_12323 ? _GEN_4 : mem_1858;
  assign _GEN_10057 = 11'h743 == _T_12323 ? _GEN_4 : mem_1859;
  assign _GEN_10058 = 11'h744 == _T_12323 ? _GEN_4 : mem_1860;
  assign _GEN_10059 = 11'h745 == _T_12323 ? _GEN_4 : mem_1861;
  assign _GEN_10060 = 11'h746 == _T_12323 ? _GEN_4 : mem_1862;
  assign _GEN_10061 = 11'h747 == _T_12323 ? _GEN_4 : mem_1863;
  assign _GEN_10062 = 11'h748 == _T_12323 ? _GEN_4 : mem_1864;
  assign _GEN_10063 = 11'h749 == _T_12323 ? _GEN_4 : mem_1865;
  assign _GEN_10064 = 11'h74a == _T_12323 ? _GEN_4 : mem_1866;
  assign _GEN_10065 = 11'h74b == _T_12323 ? _GEN_4 : mem_1867;
  assign _GEN_10066 = 11'h74c == _T_12323 ? _GEN_4 : mem_1868;
  assign _GEN_10067 = 11'h74d == _T_12323 ? _GEN_4 : mem_1869;
  assign _GEN_10068 = 11'h74e == _T_12323 ? _GEN_4 : mem_1870;
  assign _GEN_10069 = 11'h74f == _T_12323 ? _GEN_4 : mem_1871;
  assign _GEN_10070 = 11'h750 == _T_12323 ? _GEN_4 : mem_1872;
  assign _GEN_10071 = 11'h751 == _T_12323 ? _GEN_4 : mem_1873;
  assign _GEN_10072 = 11'h752 == _T_12323 ? _GEN_4 : mem_1874;
  assign _GEN_10073 = 11'h753 == _T_12323 ? _GEN_4 : mem_1875;
  assign _GEN_10074 = 11'h754 == _T_12323 ? _GEN_4 : mem_1876;
  assign _GEN_10075 = 11'h755 == _T_12323 ? _GEN_4 : mem_1877;
  assign _GEN_10076 = 11'h756 == _T_12323 ? _GEN_4 : mem_1878;
  assign _GEN_10077 = 11'h757 == _T_12323 ? _GEN_4 : mem_1879;
  assign _GEN_10078 = 11'h758 == _T_12323 ? _GEN_4 : mem_1880;
  assign _GEN_10079 = 11'h759 == _T_12323 ? _GEN_4 : mem_1881;
  assign _GEN_10080 = 11'h75a == _T_12323 ? _GEN_4 : mem_1882;
  assign _GEN_10081 = 11'h75b == _T_12323 ? _GEN_4 : mem_1883;
  assign _GEN_10082 = 11'h75c == _T_12323 ? _GEN_4 : mem_1884;
  assign _GEN_10083 = 11'h75d == _T_12323 ? _GEN_4 : mem_1885;
  assign _GEN_10084 = 11'h75e == _T_12323 ? _GEN_4 : mem_1886;
  assign _GEN_10085 = 11'h75f == _T_12323 ? _GEN_4 : mem_1887;
  assign _GEN_10086 = 11'h760 == _T_12323 ? _GEN_4 : mem_1888;
  assign _GEN_10087 = 11'h761 == _T_12323 ? _GEN_4 : mem_1889;
  assign _GEN_10088 = 11'h762 == _T_12323 ? _GEN_4 : mem_1890;
  assign _GEN_10089 = 11'h763 == _T_12323 ? _GEN_4 : mem_1891;
  assign _GEN_10090 = 11'h764 == _T_12323 ? _GEN_4 : mem_1892;
  assign _GEN_10091 = 11'h765 == _T_12323 ? _GEN_4 : mem_1893;
  assign _GEN_10092 = 11'h766 == _T_12323 ? _GEN_4 : mem_1894;
  assign _GEN_10093 = 11'h767 == _T_12323 ? _GEN_4 : mem_1895;
  assign _GEN_10094 = 11'h768 == _T_12323 ? _GEN_4 : mem_1896;
  assign _GEN_10095 = 11'h769 == _T_12323 ? _GEN_4 : mem_1897;
  assign _GEN_10096 = 11'h76a == _T_12323 ? _GEN_4 : mem_1898;
  assign _GEN_10097 = 11'h76b == _T_12323 ? _GEN_4 : mem_1899;
  assign _GEN_10098 = 11'h76c == _T_12323 ? _GEN_4 : mem_1900;
  assign _GEN_10099 = 11'h76d == _T_12323 ? _GEN_4 : mem_1901;
  assign _GEN_10100 = 11'h76e == _T_12323 ? _GEN_4 : mem_1902;
  assign _GEN_10101 = 11'h76f == _T_12323 ? _GEN_4 : mem_1903;
  assign _GEN_10102 = 11'h770 == _T_12323 ? _GEN_4 : mem_1904;
  assign _GEN_10103 = 11'h771 == _T_12323 ? _GEN_4 : mem_1905;
  assign _GEN_10104 = 11'h772 == _T_12323 ? _GEN_4 : mem_1906;
  assign _GEN_10105 = 11'h773 == _T_12323 ? _GEN_4 : mem_1907;
  assign _GEN_10106 = 11'h774 == _T_12323 ? _GEN_4 : mem_1908;
  assign _GEN_10107 = 11'h775 == _T_12323 ? _GEN_4 : mem_1909;
  assign _GEN_10108 = 11'h776 == _T_12323 ? _GEN_4 : mem_1910;
  assign _GEN_10109 = 11'h777 == _T_12323 ? _GEN_4 : mem_1911;
  assign _GEN_10110 = 11'h778 == _T_12323 ? _GEN_4 : mem_1912;
  assign _GEN_10111 = 11'h779 == _T_12323 ? _GEN_4 : mem_1913;
  assign _GEN_10112 = 11'h77a == _T_12323 ? _GEN_4 : mem_1914;
  assign _GEN_10113 = 11'h77b == _T_12323 ? _GEN_4 : mem_1915;
  assign _GEN_10114 = 11'h77c == _T_12323 ? _GEN_4 : mem_1916;
  assign _GEN_10115 = 11'h77d == _T_12323 ? _GEN_4 : mem_1917;
  assign _GEN_10116 = 11'h77e == _T_12323 ? _GEN_4 : mem_1918;
  assign _GEN_10117 = 11'h77f == _T_12323 ? _GEN_4 : mem_1919;
  assign _GEN_10118 = 11'h780 == _T_12323 ? _GEN_4 : mem_1920;
  assign _GEN_10119 = 11'h781 == _T_12323 ? _GEN_4 : mem_1921;
  assign _GEN_10120 = 11'h782 == _T_12323 ? _GEN_4 : mem_1922;
  assign _GEN_10121 = 11'h783 == _T_12323 ? _GEN_4 : mem_1923;
  assign _GEN_10122 = 11'h784 == _T_12323 ? _GEN_4 : mem_1924;
  assign _GEN_10123 = 11'h785 == _T_12323 ? _GEN_4 : mem_1925;
  assign _GEN_10124 = 11'h786 == _T_12323 ? _GEN_4 : mem_1926;
  assign _GEN_10125 = 11'h787 == _T_12323 ? _GEN_4 : mem_1927;
  assign _GEN_10126 = 11'h788 == _T_12323 ? _GEN_4 : mem_1928;
  assign _GEN_10127 = 11'h789 == _T_12323 ? _GEN_4 : mem_1929;
  assign _GEN_10128 = 11'h78a == _T_12323 ? _GEN_4 : mem_1930;
  assign _GEN_10129 = 11'h78b == _T_12323 ? _GEN_4 : mem_1931;
  assign _GEN_10130 = 11'h78c == _T_12323 ? _GEN_4 : mem_1932;
  assign _GEN_10131 = 11'h78d == _T_12323 ? _GEN_4 : mem_1933;
  assign _GEN_10132 = 11'h78e == _T_12323 ? _GEN_4 : mem_1934;
  assign _GEN_10133 = 11'h78f == _T_12323 ? _GEN_4 : mem_1935;
  assign _GEN_10134 = 11'h790 == _T_12323 ? _GEN_4 : mem_1936;
  assign _GEN_10135 = 11'h791 == _T_12323 ? _GEN_4 : mem_1937;
  assign _GEN_10136 = 11'h792 == _T_12323 ? _GEN_4 : mem_1938;
  assign _GEN_10137 = 11'h793 == _T_12323 ? _GEN_4 : mem_1939;
  assign _GEN_10138 = 11'h794 == _T_12323 ? _GEN_4 : mem_1940;
  assign _GEN_10139 = 11'h795 == _T_12323 ? _GEN_4 : mem_1941;
  assign _GEN_10140 = 11'h796 == _T_12323 ? _GEN_4 : mem_1942;
  assign _GEN_10141 = 11'h797 == _T_12323 ? _GEN_4 : mem_1943;
  assign _GEN_10142 = 11'h798 == _T_12323 ? _GEN_4 : mem_1944;
  assign _GEN_10143 = 11'h799 == _T_12323 ? _GEN_4 : mem_1945;
  assign _GEN_10144 = 11'h79a == _T_12323 ? _GEN_4 : mem_1946;
  assign _GEN_10145 = 11'h79b == _T_12323 ? _GEN_4 : mem_1947;
  assign _GEN_10146 = 11'h79c == _T_12323 ? _GEN_4 : mem_1948;
  assign _GEN_10147 = 11'h79d == _T_12323 ? _GEN_4 : mem_1949;
  assign _GEN_10148 = 11'h79e == _T_12323 ? _GEN_4 : mem_1950;
  assign _GEN_10149 = 11'h79f == _T_12323 ? _GEN_4 : mem_1951;
  assign _GEN_10150 = 11'h7a0 == _T_12323 ? _GEN_4 : mem_1952;
  assign _GEN_10151 = 11'h7a1 == _T_12323 ? _GEN_4 : mem_1953;
  assign _GEN_10152 = 11'h7a2 == _T_12323 ? _GEN_4 : mem_1954;
  assign _GEN_10153 = 11'h7a3 == _T_12323 ? _GEN_4 : mem_1955;
  assign _GEN_10154 = 11'h7a4 == _T_12323 ? _GEN_4 : mem_1956;
  assign _GEN_10155 = 11'h7a5 == _T_12323 ? _GEN_4 : mem_1957;
  assign _GEN_10156 = 11'h7a6 == _T_12323 ? _GEN_4 : mem_1958;
  assign _GEN_10157 = 11'h7a7 == _T_12323 ? _GEN_4 : mem_1959;
  assign _GEN_10158 = 11'h7a8 == _T_12323 ? _GEN_4 : mem_1960;
  assign _GEN_10159 = 11'h7a9 == _T_12323 ? _GEN_4 : mem_1961;
  assign _GEN_10160 = 11'h7aa == _T_12323 ? _GEN_4 : mem_1962;
  assign _GEN_10161 = 11'h7ab == _T_12323 ? _GEN_4 : mem_1963;
  assign _GEN_10162 = 11'h7ac == _T_12323 ? _GEN_4 : mem_1964;
  assign _GEN_10163 = 11'h7ad == _T_12323 ? _GEN_4 : mem_1965;
  assign _GEN_10164 = 11'h7ae == _T_12323 ? _GEN_4 : mem_1966;
  assign _GEN_10165 = 11'h7af == _T_12323 ? _GEN_4 : mem_1967;
  assign _GEN_10166 = 11'h7b0 == _T_12323 ? _GEN_4 : mem_1968;
  assign _GEN_10167 = 11'h7b1 == _T_12323 ? _GEN_4 : mem_1969;
  assign _GEN_10168 = 11'h7b2 == _T_12323 ? _GEN_4 : mem_1970;
  assign _GEN_10169 = 11'h7b3 == _T_12323 ? _GEN_4 : mem_1971;
  assign _GEN_10170 = 11'h7b4 == _T_12323 ? _GEN_4 : mem_1972;
  assign _GEN_10171 = 11'h7b5 == _T_12323 ? _GEN_4 : mem_1973;
  assign _GEN_10172 = 11'h7b6 == _T_12323 ? _GEN_4 : mem_1974;
  assign _GEN_10173 = 11'h7b7 == _T_12323 ? _GEN_4 : mem_1975;
  assign _GEN_10174 = 11'h7b8 == _T_12323 ? _GEN_4 : mem_1976;
  assign _GEN_10175 = 11'h7b9 == _T_12323 ? _GEN_4 : mem_1977;
  assign _GEN_10176 = 11'h7ba == _T_12323 ? _GEN_4 : mem_1978;
  assign _GEN_10177 = 11'h7bb == _T_12323 ? _GEN_4 : mem_1979;
  assign _GEN_10178 = 11'h7bc == _T_12323 ? _GEN_4 : mem_1980;
  assign _GEN_10179 = 11'h7bd == _T_12323 ? _GEN_4 : mem_1981;
  assign _GEN_10180 = 11'h7be == _T_12323 ? _GEN_4 : mem_1982;
  assign _GEN_10181 = 11'h7bf == _T_12323 ? _GEN_4 : mem_1983;
  assign _GEN_10182 = 11'h7c0 == _T_12323 ? _GEN_4 : mem_1984;
  assign _GEN_10183 = 11'h7c1 == _T_12323 ? _GEN_4 : mem_1985;
  assign _GEN_10184 = 11'h7c2 == _T_12323 ? _GEN_4 : mem_1986;
  assign _GEN_10185 = 11'h7c3 == _T_12323 ? _GEN_4 : mem_1987;
  assign _GEN_10186 = 11'h7c4 == _T_12323 ? _GEN_4 : mem_1988;
  assign _GEN_10187 = 11'h7c5 == _T_12323 ? _GEN_4 : mem_1989;
  assign _GEN_10188 = 11'h7c6 == _T_12323 ? _GEN_4 : mem_1990;
  assign _GEN_10189 = 11'h7c7 == _T_12323 ? _GEN_4 : mem_1991;
  assign _GEN_10190 = 11'h7c8 == _T_12323 ? _GEN_4 : mem_1992;
  assign _GEN_10191 = 11'h7c9 == _T_12323 ? _GEN_4 : mem_1993;
  assign _GEN_10192 = 11'h7ca == _T_12323 ? _GEN_4 : mem_1994;
  assign _GEN_10193 = 11'h7cb == _T_12323 ? _GEN_4 : mem_1995;
  assign _GEN_10194 = 11'h7cc == _T_12323 ? _GEN_4 : mem_1996;
  assign _GEN_10195 = 11'h7cd == _T_12323 ? _GEN_4 : mem_1997;
  assign _GEN_10196 = 11'h7ce == _T_12323 ? _GEN_4 : mem_1998;
  assign _GEN_10197 = 11'h7cf == _T_12323 ? _GEN_4 : mem_1999;
  assign _GEN_10198 = 11'h7d0 == _T_12323 ? _GEN_4 : mem_2000;
  assign _GEN_10199 = 11'h7d1 == _T_12323 ? _GEN_4 : mem_2001;
  assign _GEN_10200 = 11'h7d2 == _T_12323 ? _GEN_4 : mem_2002;
  assign _GEN_10201 = 11'h7d3 == _T_12323 ? _GEN_4 : mem_2003;
  assign _GEN_10202 = 11'h7d4 == _T_12323 ? _GEN_4 : mem_2004;
  assign _GEN_10203 = 11'h7d5 == _T_12323 ? _GEN_4 : mem_2005;
  assign _GEN_10204 = 11'h7d6 == _T_12323 ? _GEN_4 : mem_2006;
  assign _GEN_10205 = 11'h7d7 == _T_12323 ? _GEN_4 : mem_2007;
  assign _GEN_10206 = 11'h7d8 == _T_12323 ? _GEN_4 : mem_2008;
  assign _GEN_10207 = 11'h7d9 == _T_12323 ? _GEN_4 : mem_2009;
  assign _GEN_10208 = 11'h7da == _T_12323 ? _GEN_4 : mem_2010;
  assign _GEN_10209 = 11'h7db == _T_12323 ? _GEN_4 : mem_2011;
  assign _GEN_10210 = 11'h7dc == _T_12323 ? _GEN_4 : mem_2012;
  assign _GEN_10211 = 11'h7dd == _T_12323 ? _GEN_4 : mem_2013;
  assign _GEN_10212 = 11'h7de == _T_12323 ? _GEN_4 : mem_2014;
  assign _GEN_10213 = 11'h7df == _T_12323 ? _GEN_4 : mem_2015;
  assign _GEN_10214 = 11'h7e0 == _T_12323 ? _GEN_4 : mem_2016;
  assign _GEN_10215 = 11'h7e1 == _T_12323 ? _GEN_4 : mem_2017;
  assign _GEN_10216 = 11'h7e2 == _T_12323 ? _GEN_4 : mem_2018;
  assign _GEN_10217 = 11'h7e3 == _T_12323 ? _GEN_4 : mem_2019;
  assign _GEN_10218 = 11'h7e4 == _T_12323 ? _GEN_4 : mem_2020;
  assign _GEN_10219 = 11'h7e5 == _T_12323 ? _GEN_4 : mem_2021;
  assign _GEN_10220 = 11'h7e6 == _T_12323 ? _GEN_4 : mem_2022;
  assign _GEN_10221 = 11'h7e7 == _T_12323 ? _GEN_4 : mem_2023;
  assign _GEN_10222 = 11'h7e8 == _T_12323 ? _GEN_4 : mem_2024;
  assign _GEN_10223 = 11'h7e9 == _T_12323 ? _GEN_4 : mem_2025;
  assign _GEN_10224 = 11'h7ea == _T_12323 ? _GEN_4 : mem_2026;
  assign _GEN_10225 = 11'h7eb == _T_12323 ? _GEN_4 : mem_2027;
  assign _GEN_10226 = 11'h7ec == _T_12323 ? _GEN_4 : mem_2028;
  assign _GEN_10227 = 11'h7ed == _T_12323 ? _GEN_4 : mem_2029;
  assign _GEN_10228 = 11'h7ee == _T_12323 ? _GEN_4 : mem_2030;
  assign _GEN_10229 = 11'h7ef == _T_12323 ? _GEN_4 : mem_2031;
  assign _GEN_10230 = 11'h7f0 == _T_12323 ? _GEN_4 : mem_2032;
  assign _GEN_10231 = 11'h7f1 == _T_12323 ? _GEN_4 : mem_2033;
  assign _GEN_10232 = 11'h7f2 == _T_12323 ? _GEN_4 : mem_2034;
  assign _GEN_10233 = 11'h7f3 == _T_12323 ? _GEN_4 : mem_2035;
  assign _GEN_10234 = 11'h7f4 == _T_12323 ? _GEN_4 : mem_2036;
  assign _GEN_10235 = 11'h7f5 == _T_12323 ? _GEN_4 : mem_2037;
  assign _GEN_10236 = 11'h7f6 == _T_12323 ? _GEN_4 : mem_2038;
  assign _GEN_10237 = 11'h7f7 == _T_12323 ? _GEN_4 : mem_2039;
  assign _GEN_10238 = 11'h7f8 == _T_12323 ? _GEN_4 : mem_2040;
  assign _GEN_10239 = 11'h7f9 == _T_12323 ? _GEN_4 : mem_2041;
  assign _GEN_10240 = 11'h7fa == _T_12323 ? _GEN_4 : mem_2042;
  assign _GEN_10241 = 11'h7fb == _T_12323 ? _GEN_4 : mem_2043;
  assign _GEN_10242 = 11'h7fc == _T_12323 ? _GEN_4 : mem_2044;
  assign _GEN_10243 = 11'h7fd == _T_12323 ? _GEN_4 : mem_2045;
  assign _GEN_10244 = 11'h7fe == _T_12323 ? _GEN_4 : mem_2046;
  assign _GEN_10245 = 11'h7ff == _T_12323 ? _GEN_4 : mem_2047;
  assign rdata = _GEN_5;
  assign toWrite_0 = _GEN_2053;
  assign toWrite_1 = _GEN_4101;
  assign toWrite_2 = _GEN_6149;
  assign toWrite_3 = _GEN_8197;
  assign _GEN_0 = _GEN_2052;
  assign _GEN_1 = _GEN_2052;
  assign _GEN_2 = _GEN_2052;
  assign _GEN_3 = _GEN_2052;
  assign _GEN_4 = _T_12358;
  assign _GEN_5 = _GEN_2052;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  mem_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  mem_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  mem_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  mem_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  mem_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  mem_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  mem_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  mem_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  mem_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  mem_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  mem_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  mem_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  mem_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  mem_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  mem_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  mem_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  mem_16 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  mem_17 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  mem_18 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  mem_19 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  mem_20 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  mem_21 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  mem_22 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  mem_23 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  mem_24 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  mem_25 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  mem_26 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  mem_27 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  mem_28 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  mem_29 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  mem_30 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  mem_31 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  mem_32 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  mem_33 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  mem_34 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  mem_35 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  mem_36 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  mem_37 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  mem_38 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  mem_39 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  mem_40 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  mem_41 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  mem_42 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  mem_43 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  mem_44 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  mem_45 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  mem_46 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  mem_47 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  mem_48 = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  mem_49 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  mem_50 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  mem_51 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  mem_52 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  mem_53 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  mem_54 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  mem_55 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  mem_56 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  mem_57 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  mem_58 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  mem_59 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  mem_60 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  mem_61 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  mem_62 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  mem_63 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  mem_64 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  mem_65 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  mem_66 = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  mem_67 = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  mem_68 = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  mem_69 = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  mem_70 = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  mem_71 = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  mem_72 = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  mem_73 = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  mem_74 = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  mem_75 = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  mem_76 = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  mem_77 = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  mem_78 = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  mem_79 = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  mem_80 = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  mem_81 = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  mem_82 = _RAND_82[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  mem_83 = _RAND_83[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  mem_84 = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  mem_85 = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  mem_86 = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  mem_87 = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  mem_88 = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  mem_89 = _RAND_89[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  mem_90 = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  mem_91 = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  mem_92 = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  mem_93 = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  mem_94 = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  mem_95 = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  mem_96 = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  mem_97 = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  mem_98 = _RAND_98[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  mem_99 = _RAND_99[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  mem_100 = _RAND_100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  mem_101 = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  mem_102 = _RAND_102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  mem_103 = _RAND_103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  mem_104 = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  mem_105 = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  mem_106 = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  mem_107 = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  mem_108 = _RAND_108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  mem_109 = _RAND_109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  mem_110 = _RAND_110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  mem_111 = _RAND_111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  mem_112 = _RAND_112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  mem_113 = _RAND_113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  mem_114 = _RAND_114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  mem_115 = _RAND_115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  mem_116 = _RAND_116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  mem_117 = _RAND_117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  mem_118 = _RAND_118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  mem_119 = _RAND_119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  mem_120 = _RAND_120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  mem_121 = _RAND_121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  mem_122 = _RAND_122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  mem_123 = _RAND_123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  mem_124 = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  mem_125 = _RAND_125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  mem_126 = _RAND_126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  mem_127 = _RAND_127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  mem_128 = _RAND_128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{$random}};
  mem_129 = _RAND_129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  mem_130 = _RAND_130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{$random}};
  mem_131 = _RAND_131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{$random}};
  mem_132 = _RAND_132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{$random}};
  mem_133 = _RAND_133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{$random}};
  mem_134 = _RAND_134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{$random}};
  mem_135 = _RAND_135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{$random}};
  mem_136 = _RAND_136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{$random}};
  mem_137 = _RAND_137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{$random}};
  mem_138 = _RAND_138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{$random}};
  mem_139 = _RAND_139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{$random}};
  mem_140 = _RAND_140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{$random}};
  mem_141 = _RAND_141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{$random}};
  mem_142 = _RAND_142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{$random}};
  mem_143 = _RAND_143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{$random}};
  mem_144 = _RAND_144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{$random}};
  mem_145 = _RAND_145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{$random}};
  mem_146 = _RAND_146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{$random}};
  mem_147 = _RAND_147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{$random}};
  mem_148 = _RAND_148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{$random}};
  mem_149 = _RAND_149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{$random}};
  mem_150 = _RAND_150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{$random}};
  mem_151 = _RAND_151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{$random}};
  mem_152 = _RAND_152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{$random}};
  mem_153 = _RAND_153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{$random}};
  mem_154 = _RAND_154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{$random}};
  mem_155 = _RAND_155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{$random}};
  mem_156 = _RAND_156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{$random}};
  mem_157 = _RAND_157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{$random}};
  mem_158 = _RAND_158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{$random}};
  mem_159 = _RAND_159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{$random}};
  mem_160 = _RAND_160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{$random}};
  mem_161 = _RAND_161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{$random}};
  mem_162 = _RAND_162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{$random}};
  mem_163 = _RAND_163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{$random}};
  mem_164 = _RAND_164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{$random}};
  mem_165 = _RAND_165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{$random}};
  mem_166 = _RAND_166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{$random}};
  mem_167 = _RAND_167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{$random}};
  mem_168 = _RAND_168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{$random}};
  mem_169 = _RAND_169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{$random}};
  mem_170 = _RAND_170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{$random}};
  mem_171 = _RAND_171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{$random}};
  mem_172 = _RAND_172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{$random}};
  mem_173 = _RAND_173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{$random}};
  mem_174 = _RAND_174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{$random}};
  mem_175 = _RAND_175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{$random}};
  mem_176 = _RAND_176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{$random}};
  mem_177 = _RAND_177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{$random}};
  mem_178 = _RAND_178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{$random}};
  mem_179 = _RAND_179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{$random}};
  mem_180 = _RAND_180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{$random}};
  mem_181 = _RAND_181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{$random}};
  mem_182 = _RAND_182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{$random}};
  mem_183 = _RAND_183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{$random}};
  mem_184 = _RAND_184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{$random}};
  mem_185 = _RAND_185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{$random}};
  mem_186 = _RAND_186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{$random}};
  mem_187 = _RAND_187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{$random}};
  mem_188 = _RAND_188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{$random}};
  mem_189 = _RAND_189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{$random}};
  mem_190 = _RAND_190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{$random}};
  mem_191 = _RAND_191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{$random}};
  mem_192 = _RAND_192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{$random}};
  mem_193 = _RAND_193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{$random}};
  mem_194 = _RAND_194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{$random}};
  mem_195 = _RAND_195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{$random}};
  mem_196 = _RAND_196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{$random}};
  mem_197 = _RAND_197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{$random}};
  mem_198 = _RAND_198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{$random}};
  mem_199 = _RAND_199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{$random}};
  mem_200 = _RAND_200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{$random}};
  mem_201 = _RAND_201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{$random}};
  mem_202 = _RAND_202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{$random}};
  mem_203 = _RAND_203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{$random}};
  mem_204 = _RAND_204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{$random}};
  mem_205 = _RAND_205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{$random}};
  mem_206 = _RAND_206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{$random}};
  mem_207 = _RAND_207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{$random}};
  mem_208 = _RAND_208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{$random}};
  mem_209 = _RAND_209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{$random}};
  mem_210 = _RAND_210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{$random}};
  mem_211 = _RAND_211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{$random}};
  mem_212 = _RAND_212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{$random}};
  mem_213 = _RAND_213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{$random}};
  mem_214 = _RAND_214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{$random}};
  mem_215 = _RAND_215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{$random}};
  mem_216 = _RAND_216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{$random}};
  mem_217 = _RAND_217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{$random}};
  mem_218 = _RAND_218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{$random}};
  mem_219 = _RAND_219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{$random}};
  mem_220 = _RAND_220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{$random}};
  mem_221 = _RAND_221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{$random}};
  mem_222 = _RAND_222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{$random}};
  mem_223 = _RAND_223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{$random}};
  mem_224 = _RAND_224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{$random}};
  mem_225 = _RAND_225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{$random}};
  mem_226 = _RAND_226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{$random}};
  mem_227 = _RAND_227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{$random}};
  mem_228 = _RAND_228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{$random}};
  mem_229 = _RAND_229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{$random}};
  mem_230 = _RAND_230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{$random}};
  mem_231 = _RAND_231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{$random}};
  mem_232 = _RAND_232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{$random}};
  mem_233 = _RAND_233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{$random}};
  mem_234 = _RAND_234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{$random}};
  mem_235 = _RAND_235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{$random}};
  mem_236 = _RAND_236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{$random}};
  mem_237 = _RAND_237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{$random}};
  mem_238 = _RAND_238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{$random}};
  mem_239 = _RAND_239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{$random}};
  mem_240 = _RAND_240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{$random}};
  mem_241 = _RAND_241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{$random}};
  mem_242 = _RAND_242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{$random}};
  mem_243 = _RAND_243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{$random}};
  mem_244 = _RAND_244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{$random}};
  mem_245 = _RAND_245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{$random}};
  mem_246 = _RAND_246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{$random}};
  mem_247 = _RAND_247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{$random}};
  mem_248 = _RAND_248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{$random}};
  mem_249 = _RAND_249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{$random}};
  mem_250 = _RAND_250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{$random}};
  mem_251 = _RAND_251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{$random}};
  mem_252 = _RAND_252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{$random}};
  mem_253 = _RAND_253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{$random}};
  mem_254 = _RAND_254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{$random}};
  mem_255 = _RAND_255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{$random}};
  mem_256 = _RAND_256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{$random}};
  mem_257 = _RAND_257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{$random}};
  mem_258 = _RAND_258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{$random}};
  mem_259 = _RAND_259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{$random}};
  mem_260 = _RAND_260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{$random}};
  mem_261 = _RAND_261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{$random}};
  mem_262 = _RAND_262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{$random}};
  mem_263 = _RAND_263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{$random}};
  mem_264 = _RAND_264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{$random}};
  mem_265 = _RAND_265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{$random}};
  mem_266 = _RAND_266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{$random}};
  mem_267 = _RAND_267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{$random}};
  mem_268 = _RAND_268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{$random}};
  mem_269 = _RAND_269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{$random}};
  mem_270 = _RAND_270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{$random}};
  mem_271 = _RAND_271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{$random}};
  mem_272 = _RAND_272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{$random}};
  mem_273 = _RAND_273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{$random}};
  mem_274 = _RAND_274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{$random}};
  mem_275 = _RAND_275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{$random}};
  mem_276 = _RAND_276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{$random}};
  mem_277 = _RAND_277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{$random}};
  mem_278 = _RAND_278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{$random}};
  mem_279 = _RAND_279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{$random}};
  mem_280 = _RAND_280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{$random}};
  mem_281 = _RAND_281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{$random}};
  mem_282 = _RAND_282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{$random}};
  mem_283 = _RAND_283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{$random}};
  mem_284 = _RAND_284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{$random}};
  mem_285 = _RAND_285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{$random}};
  mem_286 = _RAND_286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{$random}};
  mem_287 = _RAND_287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{$random}};
  mem_288 = _RAND_288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{$random}};
  mem_289 = _RAND_289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{$random}};
  mem_290 = _RAND_290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{$random}};
  mem_291 = _RAND_291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{$random}};
  mem_292 = _RAND_292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{$random}};
  mem_293 = _RAND_293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{$random}};
  mem_294 = _RAND_294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{$random}};
  mem_295 = _RAND_295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{$random}};
  mem_296 = _RAND_296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{$random}};
  mem_297 = _RAND_297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{$random}};
  mem_298 = _RAND_298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{$random}};
  mem_299 = _RAND_299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{$random}};
  mem_300 = _RAND_300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{$random}};
  mem_301 = _RAND_301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{$random}};
  mem_302 = _RAND_302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{$random}};
  mem_303 = _RAND_303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{$random}};
  mem_304 = _RAND_304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{$random}};
  mem_305 = _RAND_305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{$random}};
  mem_306 = _RAND_306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{$random}};
  mem_307 = _RAND_307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{$random}};
  mem_308 = _RAND_308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{$random}};
  mem_309 = _RAND_309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{$random}};
  mem_310 = _RAND_310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{$random}};
  mem_311 = _RAND_311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{$random}};
  mem_312 = _RAND_312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{$random}};
  mem_313 = _RAND_313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{$random}};
  mem_314 = _RAND_314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{$random}};
  mem_315 = _RAND_315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{$random}};
  mem_316 = _RAND_316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{$random}};
  mem_317 = _RAND_317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{$random}};
  mem_318 = _RAND_318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{$random}};
  mem_319 = _RAND_319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{$random}};
  mem_320 = _RAND_320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{$random}};
  mem_321 = _RAND_321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{$random}};
  mem_322 = _RAND_322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{$random}};
  mem_323 = _RAND_323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{$random}};
  mem_324 = _RAND_324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{$random}};
  mem_325 = _RAND_325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{$random}};
  mem_326 = _RAND_326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{$random}};
  mem_327 = _RAND_327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{$random}};
  mem_328 = _RAND_328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{$random}};
  mem_329 = _RAND_329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{$random}};
  mem_330 = _RAND_330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{$random}};
  mem_331 = _RAND_331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{$random}};
  mem_332 = _RAND_332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{$random}};
  mem_333 = _RAND_333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{$random}};
  mem_334 = _RAND_334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{$random}};
  mem_335 = _RAND_335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{$random}};
  mem_336 = _RAND_336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{$random}};
  mem_337 = _RAND_337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{$random}};
  mem_338 = _RAND_338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{$random}};
  mem_339 = _RAND_339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{$random}};
  mem_340 = _RAND_340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{$random}};
  mem_341 = _RAND_341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{$random}};
  mem_342 = _RAND_342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{$random}};
  mem_343 = _RAND_343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{$random}};
  mem_344 = _RAND_344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{$random}};
  mem_345 = _RAND_345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{$random}};
  mem_346 = _RAND_346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{$random}};
  mem_347 = _RAND_347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{$random}};
  mem_348 = _RAND_348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{$random}};
  mem_349 = _RAND_349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{$random}};
  mem_350 = _RAND_350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{$random}};
  mem_351 = _RAND_351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{$random}};
  mem_352 = _RAND_352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{$random}};
  mem_353 = _RAND_353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{$random}};
  mem_354 = _RAND_354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{$random}};
  mem_355 = _RAND_355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{$random}};
  mem_356 = _RAND_356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{$random}};
  mem_357 = _RAND_357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{$random}};
  mem_358 = _RAND_358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{$random}};
  mem_359 = _RAND_359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{$random}};
  mem_360 = _RAND_360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{$random}};
  mem_361 = _RAND_361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{$random}};
  mem_362 = _RAND_362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{$random}};
  mem_363 = _RAND_363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{$random}};
  mem_364 = _RAND_364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{$random}};
  mem_365 = _RAND_365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{$random}};
  mem_366 = _RAND_366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{$random}};
  mem_367 = _RAND_367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{$random}};
  mem_368 = _RAND_368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{$random}};
  mem_369 = _RAND_369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{$random}};
  mem_370 = _RAND_370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{$random}};
  mem_371 = _RAND_371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{$random}};
  mem_372 = _RAND_372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{$random}};
  mem_373 = _RAND_373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{$random}};
  mem_374 = _RAND_374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{$random}};
  mem_375 = _RAND_375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{$random}};
  mem_376 = _RAND_376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{$random}};
  mem_377 = _RAND_377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{$random}};
  mem_378 = _RAND_378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{$random}};
  mem_379 = _RAND_379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{$random}};
  mem_380 = _RAND_380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{$random}};
  mem_381 = _RAND_381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{$random}};
  mem_382 = _RAND_382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{$random}};
  mem_383 = _RAND_383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{$random}};
  mem_384 = _RAND_384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{$random}};
  mem_385 = _RAND_385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{$random}};
  mem_386 = _RAND_386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{$random}};
  mem_387 = _RAND_387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{$random}};
  mem_388 = _RAND_388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{$random}};
  mem_389 = _RAND_389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{$random}};
  mem_390 = _RAND_390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{$random}};
  mem_391 = _RAND_391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{$random}};
  mem_392 = _RAND_392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{$random}};
  mem_393 = _RAND_393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{$random}};
  mem_394 = _RAND_394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{$random}};
  mem_395 = _RAND_395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{$random}};
  mem_396 = _RAND_396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{$random}};
  mem_397 = _RAND_397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{$random}};
  mem_398 = _RAND_398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{$random}};
  mem_399 = _RAND_399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{$random}};
  mem_400 = _RAND_400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{$random}};
  mem_401 = _RAND_401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{$random}};
  mem_402 = _RAND_402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{$random}};
  mem_403 = _RAND_403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{$random}};
  mem_404 = _RAND_404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{$random}};
  mem_405 = _RAND_405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{$random}};
  mem_406 = _RAND_406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{$random}};
  mem_407 = _RAND_407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{$random}};
  mem_408 = _RAND_408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{$random}};
  mem_409 = _RAND_409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{$random}};
  mem_410 = _RAND_410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{$random}};
  mem_411 = _RAND_411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{$random}};
  mem_412 = _RAND_412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{$random}};
  mem_413 = _RAND_413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{$random}};
  mem_414 = _RAND_414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{$random}};
  mem_415 = _RAND_415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{$random}};
  mem_416 = _RAND_416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{$random}};
  mem_417 = _RAND_417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{$random}};
  mem_418 = _RAND_418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{$random}};
  mem_419 = _RAND_419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{$random}};
  mem_420 = _RAND_420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{$random}};
  mem_421 = _RAND_421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{$random}};
  mem_422 = _RAND_422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{$random}};
  mem_423 = _RAND_423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{$random}};
  mem_424 = _RAND_424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{$random}};
  mem_425 = _RAND_425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{$random}};
  mem_426 = _RAND_426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{$random}};
  mem_427 = _RAND_427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{$random}};
  mem_428 = _RAND_428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{$random}};
  mem_429 = _RAND_429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{$random}};
  mem_430 = _RAND_430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{$random}};
  mem_431 = _RAND_431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{$random}};
  mem_432 = _RAND_432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{$random}};
  mem_433 = _RAND_433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{$random}};
  mem_434 = _RAND_434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{$random}};
  mem_435 = _RAND_435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{$random}};
  mem_436 = _RAND_436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{$random}};
  mem_437 = _RAND_437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{$random}};
  mem_438 = _RAND_438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{$random}};
  mem_439 = _RAND_439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{$random}};
  mem_440 = _RAND_440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{$random}};
  mem_441 = _RAND_441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{$random}};
  mem_442 = _RAND_442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{$random}};
  mem_443 = _RAND_443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{$random}};
  mem_444 = _RAND_444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{$random}};
  mem_445 = _RAND_445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{$random}};
  mem_446 = _RAND_446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{$random}};
  mem_447 = _RAND_447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{$random}};
  mem_448 = _RAND_448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{$random}};
  mem_449 = _RAND_449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{$random}};
  mem_450 = _RAND_450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{$random}};
  mem_451 = _RAND_451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{$random}};
  mem_452 = _RAND_452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{$random}};
  mem_453 = _RAND_453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{$random}};
  mem_454 = _RAND_454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{$random}};
  mem_455 = _RAND_455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{$random}};
  mem_456 = _RAND_456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{$random}};
  mem_457 = _RAND_457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{$random}};
  mem_458 = _RAND_458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{$random}};
  mem_459 = _RAND_459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{$random}};
  mem_460 = _RAND_460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{$random}};
  mem_461 = _RAND_461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{$random}};
  mem_462 = _RAND_462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{$random}};
  mem_463 = _RAND_463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{$random}};
  mem_464 = _RAND_464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{$random}};
  mem_465 = _RAND_465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{$random}};
  mem_466 = _RAND_466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{$random}};
  mem_467 = _RAND_467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{$random}};
  mem_468 = _RAND_468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{$random}};
  mem_469 = _RAND_469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{$random}};
  mem_470 = _RAND_470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{$random}};
  mem_471 = _RAND_471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{$random}};
  mem_472 = _RAND_472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{$random}};
  mem_473 = _RAND_473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{$random}};
  mem_474 = _RAND_474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{$random}};
  mem_475 = _RAND_475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{$random}};
  mem_476 = _RAND_476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{$random}};
  mem_477 = _RAND_477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{$random}};
  mem_478 = _RAND_478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{$random}};
  mem_479 = _RAND_479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{$random}};
  mem_480 = _RAND_480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{$random}};
  mem_481 = _RAND_481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{$random}};
  mem_482 = _RAND_482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{$random}};
  mem_483 = _RAND_483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{$random}};
  mem_484 = _RAND_484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{$random}};
  mem_485 = _RAND_485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{$random}};
  mem_486 = _RAND_486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{$random}};
  mem_487 = _RAND_487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{$random}};
  mem_488 = _RAND_488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{$random}};
  mem_489 = _RAND_489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{$random}};
  mem_490 = _RAND_490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{$random}};
  mem_491 = _RAND_491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{$random}};
  mem_492 = _RAND_492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{$random}};
  mem_493 = _RAND_493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{$random}};
  mem_494 = _RAND_494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{$random}};
  mem_495 = _RAND_495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{$random}};
  mem_496 = _RAND_496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{$random}};
  mem_497 = _RAND_497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{$random}};
  mem_498 = _RAND_498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{$random}};
  mem_499 = _RAND_499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{$random}};
  mem_500 = _RAND_500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{$random}};
  mem_501 = _RAND_501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{$random}};
  mem_502 = _RAND_502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{$random}};
  mem_503 = _RAND_503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{$random}};
  mem_504 = _RAND_504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{$random}};
  mem_505 = _RAND_505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{$random}};
  mem_506 = _RAND_506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{$random}};
  mem_507 = _RAND_507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{$random}};
  mem_508 = _RAND_508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{$random}};
  mem_509 = _RAND_509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{$random}};
  mem_510 = _RAND_510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{$random}};
  mem_511 = _RAND_511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{$random}};
  mem_512 = _RAND_512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{$random}};
  mem_513 = _RAND_513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{$random}};
  mem_514 = _RAND_514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{$random}};
  mem_515 = _RAND_515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{$random}};
  mem_516 = _RAND_516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{$random}};
  mem_517 = _RAND_517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{$random}};
  mem_518 = _RAND_518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{$random}};
  mem_519 = _RAND_519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{$random}};
  mem_520 = _RAND_520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{$random}};
  mem_521 = _RAND_521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{$random}};
  mem_522 = _RAND_522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{$random}};
  mem_523 = _RAND_523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{$random}};
  mem_524 = _RAND_524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{$random}};
  mem_525 = _RAND_525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{$random}};
  mem_526 = _RAND_526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{$random}};
  mem_527 = _RAND_527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{$random}};
  mem_528 = _RAND_528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{$random}};
  mem_529 = _RAND_529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{$random}};
  mem_530 = _RAND_530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{$random}};
  mem_531 = _RAND_531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{$random}};
  mem_532 = _RAND_532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{$random}};
  mem_533 = _RAND_533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{$random}};
  mem_534 = _RAND_534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{$random}};
  mem_535 = _RAND_535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{$random}};
  mem_536 = _RAND_536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{$random}};
  mem_537 = _RAND_537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{$random}};
  mem_538 = _RAND_538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{$random}};
  mem_539 = _RAND_539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{$random}};
  mem_540 = _RAND_540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{$random}};
  mem_541 = _RAND_541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{$random}};
  mem_542 = _RAND_542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{$random}};
  mem_543 = _RAND_543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{$random}};
  mem_544 = _RAND_544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{$random}};
  mem_545 = _RAND_545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{$random}};
  mem_546 = _RAND_546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{$random}};
  mem_547 = _RAND_547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{$random}};
  mem_548 = _RAND_548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{$random}};
  mem_549 = _RAND_549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{$random}};
  mem_550 = _RAND_550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{$random}};
  mem_551 = _RAND_551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{$random}};
  mem_552 = _RAND_552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{$random}};
  mem_553 = _RAND_553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{$random}};
  mem_554 = _RAND_554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{$random}};
  mem_555 = _RAND_555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{$random}};
  mem_556 = _RAND_556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{$random}};
  mem_557 = _RAND_557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{$random}};
  mem_558 = _RAND_558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{$random}};
  mem_559 = _RAND_559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{$random}};
  mem_560 = _RAND_560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{$random}};
  mem_561 = _RAND_561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{$random}};
  mem_562 = _RAND_562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{$random}};
  mem_563 = _RAND_563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{$random}};
  mem_564 = _RAND_564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{$random}};
  mem_565 = _RAND_565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{$random}};
  mem_566 = _RAND_566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{$random}};
  mem_567 = _RAND_567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{$random}};
  mem_568 = _RAND_568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{$random}};
  mem_569 = _RAND_569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{$random}};
  mem_570 = _RAND_570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{$random}};
  mem_571 = _RAND_571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{$random}};
  mem_572 = _RAND_572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{$random}};
  mem_573 = _RAND_573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{$random}};
  mem_574 = _RAND_574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{$random}};
  mem_575 = _RAND_575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{$random}};
  mem_576 = _RAND_576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{$random}};
  mem_577 = _RAND_577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{$random}};
  mem_578 = _RAND_578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{$random}};
  mem_579 = _RAND_579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{$random}};
  mem_580 = _RAND_580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{$random}};
  mem_581 = _RAND_581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{$random}};
  mem_582 = _RAND_582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{$random}};
  mem_583 = _RAND_583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{$random}};
  mem_584 = _RAND_584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{$random}};
  mem_585 = _RAND_585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{$random}};
  mem_586 = _RAND_586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{$random}};
  mem_587 = _RAND_587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{$random}};
  mem_588 = _RAND_588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{$random}};
  mem_589 = _RAND_589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{$random}};
  mem_590 = _RAND_590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{$random}};
  mem_591 = _RAND_591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{$random}};
  mem_592 = _RAND_592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{$random}};
  mem_593 = _RAND_593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{$random}};
  mem_594 = _RAND_594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{$random}};
  mem_595 = _RAND_595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{$random}};
  mem_596 = _RAND_596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{$random}};
  mem_597 = _RAND_597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{$random}};
  mem_598 = _RAND_598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{$random}};
  mem_599 = _RAND_599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{$random}};
  mem_600 = _RAND_600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{$random}};
  mem_601 = _RAND_601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{$random}};
  mem_602 = _RAND_602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{$random}};
  mem_603 = _RAND_603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{$random}};
  mem_604 = _RAND_604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{$random}};
  mem_605 = _RAND_605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{$random}};
  mem_606 = _RAND_606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{$random}};
  mem_607 = _RAND_607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{$random}};
  mem_608 = _RAND_608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{$random}};
  mem_609 = _RAND_609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{$random}};
  mem_610 = _RAND_610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{$random}};
  mem_611 = _RAND_611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{$random}};
  mem_612 = _RAND_612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{$random}};
  mem_613 = _RAND_613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{$random}};
  mem_614 = _RAND_614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{$random}};
  mem_615 = _RAND_615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{$random}};
  mem_616 = _RAND_616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{$random}};
  mem_617 = _RAND_617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{$random}};
  mem_618 = _RAND_618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{$random}};
  mem_619 = _RAND_619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{$random}};
  mem_620 = _RAND_620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{$random}};
  mem_621 = _RAND_621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{$random}};
  mem_622 = _RAND_622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{$random}};
  mem_623 = _RAND_623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{$random}};
  mem_624 = _RAND_624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{$random}};
  mem_625 = _RAND_625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{$random}};
  mem_626 = _RAND_626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{$random}};
  mem_627 = _RAND_627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{$random}};
  mem_628 = _RAND_628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{$random}};
  mem_629 = _RAND_629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{$random}};
  mem_630 = _RAND_630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{$random}};
  mem_631 = _RAND_631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{$random}};
  mem_632 = _RAND_632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{$random}};
  mem_633 = _RAND_633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{$random}};
  mem_634 = _RAND_634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{$random}};
  mem_635 = _RAND_635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{$random}};
  mem_636 = _RAND_636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{$random}};
  mem_637 = _RAND_637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{$random}};
  mem_638 = _RAND_638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{$random}};
  mem_639 = _RAND_639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{$random}};
  mem_640 = _RAND_640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{$random}};
  mem_641 = _RAND_641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{$random}};
  mem_642 = _RAND_642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{$random}};
  mem_643 = _RAND_643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{$random}};
  mem_644 = _RAND_644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{$random}};
  mem_645 = _RAND_645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{$random}};
  mem_646 = _RAND_646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{$random}};
  mem_647 = _RAND_647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{$random}};
  mem_648 = _RAND_648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{$random}};
  mem_649 = _RAND_649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{$random}};
  mem_650 = _RAND_650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{$random}};
  mem_651 = _RAND_651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{$random}};
  mem_652 = _RAND_652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{$random}};
  mem_653 = _RAND_653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{$random}};
  mem_654 = _RAND_654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{$random}};
  mem_655 = _RAND_655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{$random}};
  mem_656 = _RAND_656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{$random}};
  mem_657 = _RAND_657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{$random}};
  mem_658 = _RAND_658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{$random}};
  mem_659 = _RAND_659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{$random}};
  mem_660 = _RAND_660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{$random}};
  mem_661 = _RAND_661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{$random}};
  mem_662 = _RAND_662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{$random}};
  mem_663 = _RAND_663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{$random}};
  mem_664 = _RAND_664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{$random}};
  mem_665 = _RAND_665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{$random}};
  mem_666 = _RAND_666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{$random}};
  mem_667 = _RAND_667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{$random}};
  mem_668 = _RAND_668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{$random}};
  mem_669 = _RAND_669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{$random}};
  mem_670 = _RAND_670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{$random}};
  mem_671 = _RAND_671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{$random}};
  mem_672 = _RAND_672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{$random}};
  mem_673 = _RAND_673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{$random}};
  mem_674 = _RAND_674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{$random}};
  mem_675 = _RAND_675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{$random}};
  mem_676 = _RAND_676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{$random}};
  mem_677 = _RAND_677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{$random}};
  mem_678 = _RAND_678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{$random}};
  mem_679 = _RAND_679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{$random}};
  mem_680 = _RAND_680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_681 = {1{$random}};
  mem_681 = _RAND_681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_682 = {1{$random}};
  mem_682 = _RAND_682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{$random}};
  mem_683 = _RAND_683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{$random}};
  mem_684 = _RAND_684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{$random}};
  mem_685 = _RAND_685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{$random}};
  mem_686 = _RAND_686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{$random}};
  mem_687 = _RAND_687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{$random}};
  mem_688 = _RAND_688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{$random}};
  mem_689 = _RAND_689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{$random}};
  mem_690 = _RAND_690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{$random}};
  mem_691 = _RAND_691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{$random}};
  mem_692 = _RAND_692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{$random}};
  mem_693 = _RAND_693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{$random}};
  mem_694 = _RAND_694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{$random}};
  mem_695 = _RAND_695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{$random}};
  mem_696 = _RAND_696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{$random}};
  mem_697 = _RAND_697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{$random}};
  mem_698 = _RAND_698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{$random}};
  mem_699 = _RAND_699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{$random}};
  mem_700 = _RAND_700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{$random}};
  mem_701 = _RAND_701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{$random}};
  mem_702 = _RAND_702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{$random}};
  mem_703 = _RAND_703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{$random}};
  mem_704 = _RAND_704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{$random}};
  mem_705 = _RAND_705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{$random}};
  mem_706 = _RAND_706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{$random}};
  mem_707 = _RAND_707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{$random}};
  mem_708 = _RAND_708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{$random}};
  mem_709 = _RAND_709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{$random}};
  mem_710 = _RAND_710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{$random}};
  mem_711 = _RAND_711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{$random}};
  mem_712 = _RAND_712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{$random}};
  mem_713 = _RAND_713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{$random}};
  mem_714 = _RAND_714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{$random}};
  mem_715 = _RAND_715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{$random}};
  mem_716 = _RAND_716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{$random}};
  mem_717 = _RAND_717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{$random}};
  mem_718 = _RAND_718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{$random}};
  mem_719 = _RAND_719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{$random}};
  mem_720 = _RAND_720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{$random}};
  mem_721 = _RAND_721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{$random}};
  mem_722 = _RAND_722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_723 = {1{$random}};
  mem_723 = _RAND_723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_724 = {1{$random}};
  mem_724 = _RAND_724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_725 = {1{$random}};
  mem_725 = _RAND_725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_726 = {1{$random}};
  mem_726 = _RAND_726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_727 = {1{$random}};
  mem_727 = _RAND_727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_728 = {1{$random}};
  mem_728 = _RAND_728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_729 = {1{$random}};
  mem_729 = _RAND_729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_730 = {1{$random}};
  mem_730 = _RAND_730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_731 = {1{$random}};
  mem_731 = _RAND_731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_732 = {1{$random}};
  mem_732 = _RAND_732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_733 = {1{$random}};
  mem_733 = _RAND_733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_734 = {1{$random}};
  mem_734 = _RAND_734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_735 = {1{$random}};
  mem_735 = _RAND_735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_736 = {1{$random}};
  mem_736 = _RAND_736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_737 = {1{$random}};
  mem_737 = _RAND_737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_738 = {1{$random}};
  mem_738 = _RAND_738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_739 = {1{$random}};
  mem_739 = _RAND_739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_740 = {1{$random}};
  mem_740 = _RAND_740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_741 = {1{$random}};
  mem_741 = _RAND_741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_742 = {1{$random}};
  mem_742 = _RAND_742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_743 = {1{$random}};
  mem_743 = _RAND_743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_744 = {1{$random}};
  mem_744 = _RAND_744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_745 = {1{$random}};
  mem_745 = _RAND_745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_746 = {1{$random}};
  mem_746 = _RAND_746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_747 = {1{$random}};
  mem_747 = _RAND_747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_748 = {1{$random}};
  mem_748 = _RAND_748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_749 = {1{$random}};
  mem_749 = _RAND_749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_750 = {1{$random}};
  mem_750 = _RAND_750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_751 = {1{$random}};
  mem_751 = _RAND_751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_752 = {1{$random}};
  mem_752 = _RAND_752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_753 = {1{$random}};
  mem_753 = _RAND_753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_754 = {1{$random}};
  mem_754 = _RAND_754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_755 = {1{$random}};
  mem_755 = _RAND_755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_756 = {1{$random}};
  mem_756 = _RAND_756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_757 = {1{$random}};
  mem_757 = _RAND_757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_758 = {1{$random}};
  mem_758 = _RAND_758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_759 = {1{$random}};
  mem_759 = _RAND_759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_760 = {1{$random}};
  mem_760 = _RAND_760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_761 = {1{$random}};
  mem_761 = _RAND_761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_762 = {1{$random}};
  mem_762 = _RAND_762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_763 = {1{$random}};
  mem_763 = _RAND_763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_764 = {1{$random}};
  mem_764 = _RAND_764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_765 = {1{$random}};
  mem_765 = _RAND_765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_766 = {1{$random}};
  mem_766 = _RAND_766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_767 = {1{$random}};
  mem_767 = _RAND_767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_768 = {1{$random}};
  mem_768 = _RAND_768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_769 = {1{$random}};
  mem_769 = _RAND_769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_770 = {1{$random}};
  mem_770 = _RAND_770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_771 = {1{$random}};
  mem_771 = _RAND_771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_772 = {1{$random}};
  mem_772 = _RAND_772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_773 = {1{$random}};
  mem_773 = _RAND_773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_774 = {1{$random}};
  mem_774 = _RAND_774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_775 = {1{$random}};
  mem_775 = _RAND_775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_776 = {1{$random}};
  mem_776 = _RAND_776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_777 = {1{$random}};
  mem_777 = _RAND_777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_778 = {1{$random}};
  mem_778 = _RAND_778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_779 = {1{$random}};
  mem_779 = _RAND_779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_780 = {1{$random}};
  mem_780 = _RAND_780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_781 = {1{$random}};
  mem_781 = _RAND_781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_782 = {1{$random}};
  mem_782 = _RAND_782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_783 = {1{$random}};
  mem_783 = _RAND_783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_784 = {1{$random}};
  mem_784 = _RAND_784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_785 = {1{$random}};
  mem_785 = _RAND_785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_786 = {1{$random}};
  mem_786 = _RAND_786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_787 = {1{$random}};
  mem_787 = _RAND_787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_788 = {1{$random}};
  mem_788 = _RAND_788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_789 = {1{$random}};
  mem_789 = _RAND_789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_790 = {1{$random}};
  mem_790 = _RAND_790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_791 = {1{$random}};
  mem_791 = _RAND_791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_792 = {1{$random}};
  mem_792 = _RAND_792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_793 = {1{$random}};
  mem_793 = _RAND_793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_794 = {1{$random}};
  mem_794 = _RAND_794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_795 = {1{$random}};
  mem_795 = _RAND_795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_796 = {1{$random}};
  mem_796 = _RAND_796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_797 = {1{$random}};
  mem_797 = _RAND_797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_798 = {1{$random}};
  mem_798 = _RAND_798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_799 = {1{$random}};
  mem_799 = _RAND_799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_800 = {1{$random}};
  mem_800 = _RAND_800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_801 = {1{$random}};
  mem_801 = _RAND_801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_802 = {1{$random}};
  mem_802 = _RAND_802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_803 = {1{$random}};
  mem_803 = _RAND_803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_804 = {1{$random}};
  mem_804 = _RAND_804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_805 = {1{$random}};
  mem_805 = _RAND_805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_806 = {1{$random}};
  mem_806 = _RAND_806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_807 = {1{$random}};
  mem_807 = _RAND_807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_808 = {1{$random}};
  mem_808 = _RAND_808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_809 = {1{$random}};
  mem_809 = _RAND_809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_810 = {1{$random}};
  mem_810 = _RAND_810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_811 = {1{$random}};
  mem_811 = _RAND_811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_812 = {1{$random}};
  mem_812 = _RAND_812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_813 = {1{$random}};
  mem_813 = _RAND_813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_814 = {1{$random}};
  mem_814 = _RAND_814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_815 = {1{$random}};
  mem_815 = _RAND_815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_816 = {1{$random}};
  mem_816 = _RAND_816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_817 = {1{$random}};
  mem_817 = _RAND_817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_818 = {1{$random}};
  mem_818 = _RAND_818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_819 = {1{$random}};
  mem_819 = _RAND_819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_820 = {1{$random}};
  mem_820 = _RAND_820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_821 = {1{$random}};
  mem_821 = _RAND_821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_822 = {1{$random}};
  mem_822 = _RAND_822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_823 = {1{$random}};
  mem_823 = _RAND_823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_824 = {1{$random}};
  mem_824 = _RAND_824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_825 = {1{$random}};
  mem_825 = _RAND_825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_826 = {1{$random}};
  mem_826 = _RAND_826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_827 = {1{$random}};
  mem_827 = _RAND_827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_828 = {1{$random}};
  mem_828 = _RAND_828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_829 = {1{$random}};
  mem_829 = _RAND_829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_830 = {1{$random}};
  mem_830 = _RAND_830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_831 = {1{$random}};
  mem_831 = _RAND_831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_832 = {1{$random}};
  mem_832 = _RAND_832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_833 = {1{$random}};
  mem_833 = _RAND_833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_834 = {1{$random}};
  mem_834 = _RAND_834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_835 = {1{$random}};
  mem_835 = _RAND_835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_836 = {1{$random}};
  mem_836 = _RAND_836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_837 = {1{$random}};
  mem_837 = _RAND_837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_838 = {1{$random}};
  mem_838 = _RAND_838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_839 = {1{$random}};
  mem_839 = _RAND_839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_840 = {1{$random}};
  mem_840 = _RAND_840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_841 = {1{$random}};
  mem_841 = _RAND_841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_842 = {1{$random}};
  mem_842 = _RAND_842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_843 = {1{$random}};
  mem_843 = _RAND_843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_844 = {1{$random}};
  mem_844 = _RAND_844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_845 = {1{$random}};
  mem_845 = _RAND_845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_846 = {1{$random}};
  mem_846 = _RAND_846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_847 = {1{$random}};
  mem_847 = _RAND_847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_848 = {1{$random}};
  mem_848 = _RAND_848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_849 = {1{$random}};
  mem_849 = _RAND_849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_850 = {1{$random}};
  mem_850 = _RAND_850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_851 = {1{$random}};
  mem_851 = _RAND_851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_852 = {1{$random}};
  mem_852 = _RAND_852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_853 = {1{$random}};
  mem_853 = _RAND_853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_854 = {1{$random}};
  mem_854 = _RAND_854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_855 = {1{$random}};
  mem_855 = _RAND_855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_856 = {1{$random}};
  mem_856 = _RAND_856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_857 = {1{$random}};
  mem_857 = _RAND_857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_858 = {1{$random}};
  mem_858 = _RAND_858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_859 = {1{$random}};
  mem_859 = _RAND_859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_860 = {1{$random}};
  mem_860 = _RAND_860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_861 = {1{$random}};
  mem_861 = _RAND_861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_862 = {1{$random}};
  mem_862 = _RAND_862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_863 = {1{$random}};
  mem_863 = _RAND_863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_864 = {1{$random}};
  mem_864 = _RAND_864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_865 = {1{$random}};
  mem_865 = _RAND_865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_866 = {1{$random}};
  mem_866 = _RAND_866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_867 = {1{$random}};
  mem_867 = _RAND_867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_868 = {1{$random}};
  mem_868 = _RAND_868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_869 = {1{$random}};
  mem_869 = _RAND_869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_870 = {1{$random}};
  mem_870 = _RAND_870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_871 = {1{$random}};
  mem_871 = _RAND_871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_872 = {1{$random}};
  mem_872 = _RAND_872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_873 = {1{$random}};
  mem_873 = _RAND_873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_874 = {1{$random}};
  mem_874 = _RAND_874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_875 = {1{$random}};
  mem_875 = _RAND_875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_876 = {1{$random}};
  mem_876 = _RAND_876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_877 = {1{$random}};
  mem_877 = _RAND_877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_878 = {1{$random}};
  mem_878 = _RAND_878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_879 = {1{$random}};
  mem_879 = _RAND_879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_880 = {1{$random}};
  mem_880 = _RAND_880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_881 = {1{$random}};
  mem_881 = _RAND_881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_882 = {1{$random}};
  mem_882 = _RAND_882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_883 = {1{$random}};
  mem_883 = _RAND_883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_884 = {1{$random}};
  mem_884 = _RAND_884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_885 = {1{$random}};
  mem_885 = _RAND_885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_886 = {1{$random}};
  mem_886 = _RAND_886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_887 = {1{$random}};
  mem_887 = _RAND_887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_888 = {1{$random}};
  mem_888 = _RAND_888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_889 = {1{$random}};
  mem_889 = _RAND_889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_890 = {1{$random}};
  mem_890 = _RAND_890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_891 = {1{$random}};
  mem_891 = _RAND_891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_892 = {1{$random}};
  mem_892 = _RAND_892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_893 = {1{$random}};
  mem_893 = _RAND_893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_894 = {1{$random}};
  mem_894 = _RAND_894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_895 = {1{$random}};
  mem_895 = _RAND_895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_896 = {1{$random}};
  mem_896 = _RAND_896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_897 = {1{$random}};
  mem_897 = _RAND_897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_898 = {1{$random}};
  mem_898 = _RAND_898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_899 = {1{$random}};
  mem_899 = _RAND_899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_900 = {1{$random}};
  mem_900 = _RAND_900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_901 = {1{$random}};
  mem_901 = _RAND_901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_902 = {1{$random}};
  mem_902 = _RAND_902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_903 = {1{$random}};
  mem_903 = _RAND_903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_904 = {1{$random}};
  mem_904 = _RAND_904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_905 = {1{$random}};
  mem_905 = _RAND_905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_906 = {1{$random}};
  mem_906 = _RAND_906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_907 = {1{$random}};
  mem_907 = _RAND_907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_908 = {1{$random}};
  mem_908 = _RAND_908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_909 = {1{$random}};
  mem_909 = _RAND_909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_910 = {1{$random}};
  mem_910 = _RAND_910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_911 = {1{$random}};
  mem_911 = _RAND_911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_912 = {1{$random}};
  mem_912 = _RAND_912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_913 = {1{$random}};
  mem_913 = _RAND_913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_914 = {1{$random}};
  mem_914 = _RAND_914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_915 = {1{$random}};
  mem_915 = _RAND_915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_916 = {1{$random}};
  mem_916 = _RAND_916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_917 = {1{$random}};
  mem_917 = _RAND_917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_918 = {1{$random}};
  mem_918 = _RAND_918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_919 = {1{$random}};
  mem_919 = _RAND_919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_920 = {1{$random}};
  mem_920 = _RAND_920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_921 = {1{$random}};
  mem_921 = _RAND_921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_922 = {1{$random}};
  mem_922 = _RAND_922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_923 = {1{$random}};
  mem_923 = _RAND_923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_924 = {1{$random}};
  mem_924 = _RAND_924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_925 = {1{$random}};
  mem_925 = _RAND_925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_926 = {1{$random}};
  mem_926 = _RAND_926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_927 = {1{$random}};
  mem_927 = _RAND_927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_928 = {1{$random}};
  mem_928 = _RAND_928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_929 = {1{$random}};
  mem_929 = _RAND_929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_930 = {1{$random}};
  mem_930 = _RAND_930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_931 = {1{$random}};
  mem_931 = _RAND_931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_932 = {1{$random}};
  mem_932 = _RAND_932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_933 = {1{$random}};
  mem_933 = _RAND_933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_934 = {1{$random}};
  mem_934 = _RAND_934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_935 = {1{$random}};
  mem_935 = _RAND_935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_936 = {1{$random}};
  mem_936 = _RAND_936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_937 = {1{$random}};
  mem_937 = _RAND_937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_938 = {1{$random}};
  mem_938 = _RAND_938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_939 = {1{$random}};
  mem_939 = _RAND_939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_940 = {1{$random}};
  mem_940 = _RAND_940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_941 = {1{$random}};
  mem_941 = _RAND_941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_942 = {1{$random}};
  mem_942 = _RAND_942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_943 = {1{$random}};
  mem_943 = _RAND_943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_944 = {1{$random}};
  mem_944 = _RAND_944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_945 = {1{$random}};
  mem_945 = _RAND_945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_946 = {1{$random}};
  mem_946 = _RAND_946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_947 = {1{$random}};
  mem_947 = _RAND_947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_948 = {1{$random}};
  mem_948 = _RAND_948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_949 = {1{$random}};
  mem_949 = _RAND_949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_950 = {1{$random}};
  mem_950 = _RAND_950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_951 = {1{$random}};
  mem_951 = _RAND_951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_952 = {1{$random}};
  mem_952 = _RAND_952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_953 = {1{$random}};
  mem_953 = _RAND_953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_954 = {1{$random}};
  mem_954 = _RAND_954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_955 = {1{$random}};
  mem_955 = _RAND_955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_956 = {1{$random}};
  mem_956 = _RAND_956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_957 = {1{$random}};
  mem_957 = _RAND_957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_958 = {1{$random}};
  mem_958 = _RAND_958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_959 = {1{$random}};
  mem_959 = _RAND_959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_960 = {1{$random}};
  mem_960 = _RAND_960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_961 = {1{$random}};
  mem_961 = _RAND_961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_962 = {1{$random}};
  mem_962 = _RAND_962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_963 = {1{$random}};
  mem_963 = _RAND_963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_964 = {1{$random}};
  mem_964 = _RAND_964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_965 = {1{$random}};
  mem_965 = _RAND_965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_966 = {1{$random}};
  mem_966 = _RAND_966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_967 = {1{$random}};
  mem_967 = _RAND_967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_968 = {1{$random}};
  mem_968 = _RAND_968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_969 = {1{$random}};
  mem_969 = _RAND_969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_970 = {1{$random}};
  mem_970 = _RAND_970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_971 = {1{$random}};
  mem_971 = _RAND_971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_972 = {1{$random}};
  mem_972 = _RAND_972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_973 = {1{$random}};
  mem_973 = _RAND_973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_974 = {1{$random}};
  mem_974 = _RAND_974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_975 = {1{$random}};
  mem_975 = _RAND_975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_976 = {1{$random}};
  mem_976 = _RAND_976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_977 = {1{$random}};
  mem_977 = _RAND_977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_978 = {1{$random}};
  mem_978 = _RAND_978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_979 = {1{$random}};
  mem_979 = _RAND_979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_980 = {1{$random}};
  mem_980 = _RAND_980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_981 = {1{$random}};
  mem_981 = _RAND_981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_982 = {1{$random}};
  mem_982 = _RAND_982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_983 = {1{$random}};
  mem_983 = _RAND_983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_984 = {1{$random}};
  mem_984 = _RAND_984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_985 = {1{$random}};
  mem_985 = _RAND_985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_986 = {1{$random}};
  mem_986 = _RAND_986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_987 = {1{$random}};
  mem_987 = _RAND_987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_988 = {1{$random}};
  mem_988 = _RAND_988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_989 = {1{$random}};
  mem_989 = _RAND_989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_990 = {1{$random}};
  mem_990 = _RAND_990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_991 = {1{$random}};
  mem_991 = _RAND_991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_992 = {1{$random}};
  mem_992 = _RAND_992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_993 = {1{$random}};
  mem_993 = _RAND_993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_994 = {1{$random}};
  mem_994 = _RAND_994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_995 = {1{$random}};
  mem_995 = _RAND_995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_996 = {1{$random}};
  mem_996 = _RAND_996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_997 = {1{$random}};
  mem_997 = _RAND_997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_998 = {1{$random}};
  mem_998 = _RAND_998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_999 = {1{$random}};
  mem_999 = _RAND_999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1000 = {1{$random}};
  mem_1000 = _RAND_1000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1001 = {1{$random}};
  mem_1001 = _RAND_1001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1002 = {1{$random}};
  mem_1002 = _RAND_1002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1003 = {1{$random}};
  mem_1003 = _RAND_1003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1004 = {1{$random}};
  mem_1004 = _RAND_1004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1005 = {1{$random}};
  mem_1005 = _RAND_1005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1006 = {1{$random}};
  mem_1006 = _RAND_1006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1007 = {1{$random}};
  mem_1007 = _RAND_1007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1008 = {1{$random}};
  mem_1008 = _RAND_1008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1009 = {1{$random}};
  mem_1009 = _RAND_1009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1010 = {1{$random}};
  mem_1010 = _RAND_1010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1011 = {1{$random}};
  mem_1011 = _RAND_1011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1012 = {1{$random}};
  mem_1012 = _RAND_1012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1013 = {1{$random}};
  mem_1013 = _RAND_1013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1014 = {1{$random}};
  mem_1014 = _RAND_1014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1015 = {1{$random}};
  mem_1015 = _RAND_1015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1016 = {1{$random}};
  mem_1016 = _RAND_1016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1017 = {1{$random}};
  mem_1017 = _RAND_1017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1018 = {1{$random}};
  mem_1018 = _RAND_1018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1019 = {1{$random}};
  mem_1019 = _RAND_1019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1020 = {1{$random}};
  mem_1020 = _RAND_1020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1021 = {1{$random}};
  mem_1021 = _RAND_1021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1022 = {1{$random}};
  mem_1022 = _RAND_1022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1023 = {1{$random}};
  mem_1023 = _RAND_1023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1024 = {1{$random}};
  mem_1024 = _RAND_1024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1025 = {1{$random}};
  mem_1025 = _RAND_1025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1026 = {1{$random}};
  mem_1026 = _RAND_1026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1027 = {1{$random}};
  mem_1027 = _RAND_1027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1028 = {1{$random}};
  mem_1028 = _RAND_1028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1029 = {1{$random}};
  mem_1029 = _RAND_1029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1030 = {1{$random}};
  mem_1030 = _RAND_1030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1031 = {1{$random}};
  mem_1031 = _RAND_1031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1032 = {1{$random}};
  mem_1032 = _RAND_1032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1033 = {1{$random}};
  mem_1033 = _RAND_1033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1034 = {1{$random}};
  mem_1034 = _RAND_1034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1035 = {1{$random}};
  mem_1035 = _RAND_1035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1036 = {1{$random}};
  mem_1036 = _RAND_1036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1037 = {1{$random}};
  mem_1037 = _RAND_1037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1038 = {1{$random}};
  mem_1038 = _RAND_1038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1039 = {1{$random}};
  mem_1039 = _RAND_1039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1040 = {1{$random}};
  mem_1040 = _RAND_1040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1041 = {1{$random}};
  mem_1041 = _RAND_1041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1042 = {1{$random}};
  mem_1042 = _RAND_1042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1043 = {1{$random}};
  mem_1043 = _RAND_1043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1044 = {1{$random}};
  mem_1044 = _RAND_1044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1045 = {1{$random}};
  mem_1045 = _RAND_1045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1046 = {1{$random}};
  mem_1046 = _RAND_1046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1047 = {1{$random}};
  mem_1047 = _RAND_1047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1048 = {1{$random}};
  mem_1048 = _RAND_1048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1049 = {1{$random}};
  mem_1049 = _RAND_1049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1050 = {1{$random}};
  mem_1050 = _RAND_1050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1051 = {1{$random}};
  mem_1051 = _RAND_1051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1052 = {1{$random}};
  mem_1052 = _RAND_1052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1053 = {1{$random}};
  mem_1053 = _RAND_1053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1054 = {1{$random}};
  mem_1054 = _RAND_1054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1055 = {1{$random}};
  mem_1055 = _RAND_1055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1056 = {1{$random}};
  mem_1056 = _RAND_1056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1057 = {1{$random}};
  mem_1057 = _RAND_1057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1058 = {1{$random}};
  mem_1058 = _RAND_1058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1059 = {1{$random}};
  mem_1059 = _RAND_1059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1060 = {1{$random}};
  mem_1060 = _RAND_1060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1061 = {1{$random}};
  mem_1061 = _RAND_1061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1062 = {1{$random}};
  mem_1062 = _RAND_1062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1063 = {1{$random}};
  mem_1063 = _RAND_1063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1064 = {1{$random}};
  mem_1064 = _RAND_1064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1065 = {1{$random}};
  mem_1065 = _RAND_1065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1066 = {1{$random}};
  mem_1066 = _RAND_1066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1067 = {1{$random}};
  mem_1067 = _RAND_1067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1068 = {1{$random}};
  mem_1068 = _RAND_1068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1069 = {1{$random}};
  mem_1069 = _RAND_1069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1070 = {1{$random}};
  mem_1070 = _RAND_1070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1071 = {1{$random}};
  mem_1071 = _RAND_1071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1072 = {1{$random}};
  mem_1072 = _RAND_1072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1073 = {1{$random}};
  mem_1073 = _RAND_1073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1074 = {1{$random}};
  mem_1074 = _RAND_1074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1075 = {1{$random}};
  mem_1075 = _RAND_1075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1076 = {1{$random}};
  mem_1076 = _RAND_1076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1077 = {1{$random}};
  mem_1077 = _RAND_1077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1078 = {1{$random}};
  mem_1078 = _RAND_1078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1079 = {1{$random}};
  mem_1079 = _RAND_1079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1080 = {1{$random}};
  mem_1080 = _RAND_1080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1081 = {1{$random}};
  mem_1081 = _RAND_1081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1082 = {1{$random}};
  mem_1082 = _RAND_1082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1083 = {1{$random}};
  mem_1083 = _RAND_1083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1084 = {1{$random}};
  mem_1084 = _RAND_1084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1085 = {1{$random}};
  mem_1085 = _RAND_1085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1086 = {1{$random}};
  mem_1086 = _RAND_1086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1087 = {1{$random}};
  mem_1087 = _RAND_1087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1088 = {1{$random}};
  mem_1088 = _RAND_1088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1089 = {1{$random}};
  mem_1089 = _RAND_1089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1090 = {1{$random}};
  mem_1090 = _RAND_1090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1091 = {1{$random}};
  mem_1091 = _RAND_1091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1092 = {1{$random}};
  mem_1092 = _RAND_1092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1093 = {1{$random}};
  mem_1093 = _RAND_1093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1094 = {1{$random}};
  mem_1094 = _RAND_1094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1095 = {1{$random}};
  mem_1095 = _RAND_1095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1096 = {1{$random}};
  mem_1096 = _RAND_1096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1097 = {1{$random}};
  mem_1097 = _RAND_1097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1098 = {1{$random}};
  mem_1098 = _RAND_1098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1099 = {1{$random}};
  mem_1099 = _RAND_1099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1100 = {1{$random}};
  mem_1100 = _RAND_1100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1101 = {1{$random}};
  mem_1101 = _RAND_1101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1102 = {1{$random}};
  mem_1102 = _RAND_1102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1103 = {1{$random}};
  mem_1103 = _RAND_1103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1104 = {1{$random}};
  mem_1104 = _RAND_1104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1105 = {1{$random}};
  mem_1105 = _RAND_1105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1106 = {1{$random}};
  mem_1106 = _RAND_1106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1107 = {1{$random}};
  mem_1107 = _RAND_1107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1108 = {1{$random}};
  mem_1108 = _RAND_1108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1109 = {1{$random}};
  mem_1109 = _RAND_1109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1110 = {1{$random}};
  mem_1110 = _RAND_1110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1111 = {1{$random}};
  mem_1111 = _RAND_1111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1112 = {1{$random}};
  mem_1112 = _RAND_1112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1113 = {1{$random}};
  mem_1113 = _RAND_1113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1114 = {1{$random}};
  mem_1114 = _RAND_1114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1115 = {1{$random}};
  mem_1115 = _RAND_1115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1116 = {1{$random}};
  mem_1116 = _RAND_1116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1117 = {1{$random}};
  mem_1117 = _RAND_1117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1118 = {1{$random}};
  mem_1118 = _RAND_1118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1119 = {1{$random}};
  mem_1119 = _RAND_1119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1120 = {1{$random}};
  mem_1120 = _RAND_1120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1121 = {1{$random}};
  mem_1121 = _RAND_1121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1122 = {1{$random}};
  mem_1122 = _RAND_1122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1123 = {1{$random}};
  mem_1123 = _RAND_1123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1124 = {1{$random}};
  mem_1124 = _RAND_1124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1125 = {1{$random}};
  mem_1125 = _RAND_1125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1126 = {1{$random}};
  mem_1126 = _RAND_1126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1127 = {1{$random}};
  mem_1127 = _RAND_1127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1128 = {1{$random}};
  mem_1128 = _RAND_1128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1129 = {1{$random}};
  mem_1129 = _RAND_1129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1130 = {1{$random}};
  mem_1130 = _RAND_1130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1131 = {1{$random}};
  mem_1131 = _RAND_1131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1132 = {1{$random}};
  mem_1132 = _RAND_1132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1133 = {1{$random}};
  mem_1133 = _RAND_1133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1134 = {1{$random}};
  mem_1134 = _RAND_1134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1135 = {1{$random}};
  mem_1135 = _RAND_1135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1136 = {1{$random}};
  mem_1136 = _RAND_1136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1137 = {1{$random}};
  mem_1137 = _RAND_1137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1138 = {1{$random}};
  mem_1138 = _RAND_1138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1139 = {1{$random}};
  mem_1139 = _RAND_1139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1140 = {1{$random}};
  mem_1140 = _RAND_1140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1141 = {1{$random}};
  mem_1141 = _RAND_1141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1142 = {1{$random}};
  mem_1142 = _RAND_1142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1143 = {1{$random}};
  mem_1143 = _RAND_1143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1144 = {1{$random}};
  mem_1144 = _RAND_1144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1145 = {1{$random}};
  mem_1145 = _RAND_1145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1146 = {1{$random}};
  mem_1146 = _RAND_1146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1147 = {1{$random}};
  mem_1147 = _RAND_1147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1148 = {1{$random}};
  mem_1148 = _RAND_1148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1149 = {1{$random}};
  mem_1149 = _RAND_1149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1150 = {1{$random}};
  mem_1150 = _RAND_1150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1151 = {1{$random}};
  mem_1151 = _RAND_1151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1152 = {1{$random}};
  mem_1152 = _RAND_1152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1153 = {1{$random}};
  mem_1153 = _RAND_1153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1154 = {1{$random}};
  mem_1154 = _RAND_1154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1155 = {1{$random}};
  mem_1155 = _RAND_1155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1156 = {1{$random}};
  mem_1156 = _RAND_1156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1157 = {1{$random}};
  mem_1157 = _RAND_1157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1158 = {1{$random}};
  mem_1158 = _RAND_1158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1159 = {1{$random}};
  mem_1159 = _RAND_1159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1160 = {1{$random}};
  mem_1160 = _RAND_1160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1161 = {1{$random}};
  mem_1161 = _RAND_1161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1162 = {1{$random}};
  mem_1162 = _RAND_1162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1163 = {1{$random}};
  mem_1163 = _RAND_1163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1164 = {1{$random}};
  mem_1164 = _RAND_1164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1165 = {1{$random}};
  mem_1165 = _RAND_1165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1166 = {1{$random}};
  mem_1166 = _RAND_1166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1167 = {1{$random}};
  mem_1167 = _RAND_1167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1168 = {1{$random}};
  mem_1168 = _RAND_1168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1169 = {1{$random}};
  mem_1169 = _RAND_1169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1170 = {1{$random}};
  mem_1170 = _RAND_1170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1171 = {1{$random}};
  mem_1171 = _RAND_1171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1172 = {1{$random}};
  mem_1172 = _RAND_1172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1173 = {1{$random}};
  mem_1173 = _RAND_1173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1174 = {1{$random}};
  mem_1174 = _RAND_1174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1175 = {1{$random}};
  mem_1175 = _RAND_1175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1176 = {1{$random}};
  mem_1176 = _RAND_1176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1177 = {1{$random}};
  mem_1177 = _RAND_1177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1178 = {1{$random}};
  mem_1178 = _RAND_1178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1179 = {1{$random}};
  mem_1179 = _RAND_1179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1180 = {1{$random}};
  mem_1180 = _RAND_1180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1181 = {1{$random}};
  mem_1181 = _RAND_1181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1182 = {1{$random}};
  mem_1182 = _RAND_1182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1183 = {1{$random}};
  mem_1183 = _RAND_1183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1184 = {1{$random}};
  mem_1184 = _RAND_1184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1185 = {1{$random}};
  mem_1185 = _RAND_1185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1186 = {1{$random}};
  mem_1186 = _RAND_1186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1187 = {1{$random}};
  mem_1187 = _RAND_1187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1188 = {1{$random}};
  mem_1188 = _RAND_1188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1189 = {1{$random}};
  mem_1189 = _RAND_1189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1190 = {1{$random}};
  mem_1190 = _RAND_1190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1191 = {1{$random}};
  mem_1191 = _RAND_1191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1192 = {1{$random}};
  mem_1192 = _RAND_1192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1193 = {1{$random}};
  mem_1193 = _RAND_1193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1194 = {1{$random}};
  mem_1194 = _RAND_1194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1195 = {1{$random}};
  mem_1195 = _RAND_1195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1196 = {1{$random}};
  mem_1196 = _RAND_1196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1197 = {1{$random}};
  mem_1197 = _RAND_1197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1198 = {1{$random}};
  mem_1198 = _RAND_1198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1199 = {1{$random}};
  mem_1199 = _RAND_1199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1200 = {1{$random}};
  mem_1200 = _RAND_1200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1201 = {1{$random}};
  mem_1201 = _RAND_1201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1202 = {1{$random}};
  mem_1202 = _RAND_1202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1203 = {1{$random}};
  mem_1203 = _RAND_1203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1204 = {1{$random}};
  mem_1204 = _RAND_1204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1205 = {1{$random}};
  mem_1205 = _RAND_1205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1206 = {1{$random}};
  mem_1206 = _RAND_1206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1207 = {1{$random}};
  mem_1207 = _RAND_1207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1208 = {1{$random}};
  mem_1208 = _RAND_1208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1209 = {1{$random}};
  mem_1209 = _RAND_1209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1210 = {1{$random}};
  mem_1210 = _RAND_1210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1211 = {1{$random}};
  mem_1211 = _RAND_1211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1212 = {1{$random}};
  mem_1212 = _RAND_1212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1213 = {1{$random}};
  mem_1213 = _RAND_1213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1214 = {1{$random}};
  mem_1214 = _RAND_1214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1215 = {1{$random}};
  mem_1215 = _RAND_1215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1216 = {1{$random}};
  mem_1216 = _RAND_1216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1217 = {1{$random}};
  mem_1217 = _RAND_1217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1218 = {1{$random}};
  mem_1218 = _RAND_1218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1219 = {1{$random}};
  mem_1219 = _RAND_1219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1220 = {1{$random}};
  mem_1220 = _RAND_1220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1221 = {1{$random}};
  mem_1221 = _RAND_1221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1222 = {1{$random}};
  mem_1222 = _RAND_1222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1223 = {1{$random}};
  mem_1223 = _RAND_1223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1224 = {1{$random}};
  mem_1224 = _RAND_1224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1225 = {1{$random}};
  mem_1225 = _RAND_1225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1226 = {1{$random}};
  mem_1226 = _RAND_1226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1227 = {1{$random}};
  mem_1227 = _RAND_1227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1228 = {1{$random}};
  mem_1228 = _RAND_1228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1229 = {1{$random}};
  mem_1229 = _RAND_1229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1230 = {1{$random}};
  mem_1230 = _RAND_1230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1231 = {1{$random}};
  mem_1231 = _RAND_1231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1232 = {1{$random}};
  mem_1232 = _RAND_1232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1233 = {1{$random}};
  mem_1233 = _RAND_1233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1234 = {1{$random}};
  mem_1234 = _RAND_1234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1235 = {1{$random}};
  mem_1235 = _RAND_1235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1236 = {1{$random}};
  mem_1236 = _RAND_1236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1237 = {1{$random}};
  mem_1237 = _RAND_1237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1238 = {1{$random}};
  mem_1238 = _RAND_1238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1239 = {1{$random}};
  mem_1239 = _RAND_1239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1240 = {1{$random}};
  mem_1240 = _RAND_1240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1241 = {1{$random}};
  mem_1241 = _RAND_1241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1242 = {1{$random}};
  mem_1242 = _RAND_1242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1243 = {1{$random}};
  mem_1243 = _RAND_1243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1244 = {1{$random}};
  mem_1244 = _RAND_1244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1245 = {1{$random}};
  mem_1245 = _RAND_1245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1246 = {1{$random}};
  mem_1246 = _RAND_1246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1247 = {1{$random}};
  mem_1247 = _RAND_1247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1248 = {1{$random}};
  mem_1248 = _RAND_1248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1249 = {1{$random}};
  mem_1249 = _RAND_1249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1250 = {1{$random}};
  mem_1250 = _RAND_1250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1251 = {1{$random}};
  mem_1251 = _RAND_1251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1252 = {1{$random}};
  mem_1252 = _RAND_1252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1253 = {1{$random}};
  mem_1253 = _RAND_1253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1254 = {1{$random}};
  mem_1254 = _RAND_1254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1255 = {1{$random}};
  mem_1255 = _RAND_1255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1256 = {1{$random}};
  mem_1256 = _RAND_1256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1257 = {1{$random}};
  mem_1257 = _RAND_1257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1258 = {1{$random}};
  mem_1258 = _RAND_1258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1259 = {1{$random}};
  mem_1259 = _RAND_1259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1260 = {1{$random}};
  mem_1260 = _RAND_1260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1261 = {1{$random}};
  mem_1261 = _RAND_1261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1262 = {1{$random}};
  mem_1262 = _RAND_1262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1263 = {1{$random}};
  mem_1263 = _RAND_1263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1264 = {1{$random}};
  mem_1264 = _RAND_1264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1265 = {1{$random}};
  mem_1265 = _RAND_1265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1266 = {1{$random}};
  mem_1266 = _RAND_1266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1267 = {1{$random}};
  mem_1267 = _RAND_1267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1268 = {1{$random}};
  mem_1268 = _RAND_1268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1269 = {1{$random}};
  mem_1269 = _RAND_1269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1270 = {1{$random}};
  mem_1270 = _RAND_1270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1271 = {1{$random}};
  mem_1271 = _RAND_1271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1272 = {1{$random}};
  mem_1272 = _RAND_1272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1273 = {1{$random}};
  mem_1273 = _RAND_1273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1274 = {1{$random}};
  mem_1274 = _RAND_1274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1275 = {1{$random}};
  mem_1275 = _RAND_1275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1276 = {1{$random}};
  mem_1276 = _RAND_1276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1277 = {1{$random}};
  mem_1277 = _RAND_1277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1278 = {1{$random}};
  mem_1278 = _RAND_1278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1279 = {1{$random}};
  mem_1279 = _RAND_1279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1280 = {1{$random}};
  mem_1280 = _RAND_1280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1281 = {1{$random}};
  mem_1281 = _RAND_1281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1282 = {1{$random}};
  mem_1282 = _RAND_1282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1283 = {1{$random}};
  mem_1283 = _RAND_1283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1284 = {1{$random}};
  mem_1284 = _RAND_1284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1285 = {1{$random}};
  mem_1285 = _RAND_1285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1286 = {1{$random}};
  mem_1286 = _RAND_1286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1287 = {1{$random}};
  mem_1287 = _RAND_1287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1288 = {1{$random}};
  mem_1288 = _RAND_1288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1289 = {1{$random}};
  mem_1289 = _RAND_1289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1290 = {1{$random}};
  mem_1290 = _RAND_1290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1291 = {1{$random}};
  mem_1291 = _RAND_1291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1292 = {1{$random}};
  mem_1292 = _RAND_1292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1293 = {1{$random}};
  mem_1293 = _RAND_1293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1294 = {1{$random}};
  mem_1294 = _RAND_1294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1295 = {1{$random}};
  mem_1295 = _RAND_1295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1296 = {1{$random}};
  mem_1296 = _RAND_1296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1297 = {1{$random}};
  mem_1297 = _RAND_1297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1298 = {1{$random}};
  mem_1298 = _RAND_1298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1299 = {1{$random}};
  mem_1299 = _RAND_1299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1300 = {1{$random}};
  mem_1300 = _RAND_1300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1301 = {1{$random}};
  mem_1301 = _RAND_1301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1302 = {1{$random}};
  mem_1302 = _RAND_1302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1303 = {1{$random}};
  mem_1303 = _RAND_1303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1304 = {1{$random}};
  mem_1304 = _RAND_1304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1305 = {1{$random}};
  mem_1305 = _RAND_1305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1306 = {1{$random}};
  mem_1306 = _RAND_1306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1307 = {1{$random}};
  mem_1307 = _RAND_1307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1308 = {1{$random}};
  mem_1308 = _RAND_1308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1309 = {1{$random}};
  mem_1309 = _RAND_1309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1310 = {1{$random}};
  mem_1310 = _RAND_1310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1311 = {1{$random}};
  mem_1311 = _RAND_1311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1312 = {1{$random}};
  mem_1312 = _RAND_1312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1313 = {1{$random}};
  mem_1313 = _RAND_1313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1314 = {1{$random}};
  mem_1314 = _RAND_1314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1315 = {1{$random}};
  mem_1315 = _RAND_1315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1316 = {1{$random}};
  mem_1316 = _RAND_1316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1317 = {1{$random}};
  mem_1317 = _RAND_1317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1318 = {1{$random}};
  mem_1318 = _RAND_1318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1319 = {1{$random}};
  mem_1319 = _RAND_1319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1320 = {1{$random}};
  mem_1320 = _RAND_1320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1321 = {1{$random}};
  mem_1321 = _RAND_1321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1322 = {1{$random}};
  mem_1322 = _RAND_1322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1323 = {1{$random}};
  mem_1323 = _RAND_1323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1324 = {1{$random}};
  mem_1324 = _RAND_1324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1325 = {1{$random}};
  mem_1325 = _RAND_1325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1326 = {1{$random}};
  mem_1326 = _RAND_1326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1327 = {1{$random}};
  mem_1327 = _RAND_1327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1328 = {1{$random}};
  mem_1328 = _RAND_1328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1329 = {1{$random}};
  mem_1329 = _RAND_1329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1330 = {1{$random}};
  mem_1330 = _RAND_1330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1331 = {1{$random}};
  mem_1331 = _RAND_1331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1332 = {1{$random}};
  mem_1332 = _RAND_1332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1333 = {1{$random}};
  mem_1333 = _RAND_1333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1334 = {1{$random}};
  mem_1334 = _RAND_1334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1335 = {1{$random}};
  mem_1335 = _RAND_1335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1336 = {1{$random}};
  mem_1336 = _RAND_1336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1337 = {1{$random}};
  mem_1337 = _RAND_1337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1338 = {1{$random}};
  mem_1338 = _RAND_1338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1339 = {1{$random}};
  mem_1339 = _RAND_1339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1340 = {1{$random}};
  mem_1340 = _RAND_1340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1341 = {1{$random}};
  mem_1341 = _RAND_1341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1342 = {1{$random}};
  mem_1342 = _RAND_1342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1343 = {1{$random}};
  mem_1343 = _RAND_1343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1344 = {1{$random}};
  mem_1344 = _RAND_1344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1345 = {1{$random}};
  mem_1345 = _RAND_1345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1346 = {1{$random}};
  mem_1346 = _RAND_1346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1347 = {1{$random}};
  mem_1347 = _RAND_1347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1348 = {1{$random}};
  mem_1348 = _RAND_1348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1349 = {1{$random}};
  mem_1349 = _RAND_1349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1350 = {1{$random}};
  mem_1350 = _RAND_1350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1351 = {1{$random}};
  mem_1351 = _RAND_1351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1352 = {1{$random}};
  mem_1352 = _RAND_1352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1353 = {1{$random}};
  mem_1353 = _RAND_1353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1354 = {1{$random}};
  mem_1354 = _RAND_1354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1355 = {1{$random}};
  mem_1355 = _RAND_1355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1356 = {1{$random}};
  mem_1356 = _RAND_1356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1357 = {1{$random}};
  mem_1357 = _RAND_1357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1358 = {1{$random}};
  mem_1358 = _RAND_1358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1359 = {1{$random}};
  mem_1359 = _RAND_1359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1360 = {1{$random}};
  mem_1360 = _RAND_1360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1361 = {1{$random}};
  mem_1361 = _RAND_1361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1362 = {1{$random}};
  mem_1362 = _RAND_1362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1363 = {1{$random}};
  mem_1363 = _RAND_1363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1364 = {1{$random}};
  mem_1364 = _RAND_1364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1365 = {1{$random}};
  mem_1365 = _RAND_1365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1366 = {1{$random}};
  mem_1366 = _RAND_1366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1367 = {1{$random}};
  mem_1367 = _RAND_1367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1368 = {1{$random}};
  mem_1368 = _RAND_1368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1369 = {1{$random}};
  mem_1369 = _RAND_1369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1370 = {1{$random}};
  mem_1370 = _RAND_1370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1371 = {1{$random}};
  mem_1371 = _RAND_1371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1372 = {1{$random}};
  mem_1372 = _RAND_1372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1373 = {1{$random}};
  mem_1373 = _RAND_1373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1374 = {1{$random}};
  mem_1374 = _RAND_1374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1375 = {1{$random}};
  mem_1375 = _RAND_1375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1376 = {1{$random}};
  mem_1376 = _RAND_1376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1377 = {1{$random}};
  mem_1377 = _RAND_1377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1378 = {1{$random}};
  mem_1378 = _RAND_1378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1379 = {1{$random}};
  mem_1379 = _RAND_1379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1380 = {1{$random}};
  mem_1380 = _RAND_1380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1381 = {1{$random}};
  mem_1381 = _RAND_1381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1382 = {1{$random}};
  mem_1382 = _RAND_1382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1383 = {1{$random}};
  mem_1383 = _RAND_1383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1384 = {1{$random}};
  mem_1384 = _RAND_1384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1385 = {1{$random}};
  mem_1385 = _RAND_1385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1386 = {1{$random}};
  mem_1386 = _RAND_1386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1387 = {1{$random}};
  mem_1387 = _RAND_1387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1388 = {1{$random}};
  mem_1388 = _RAND_1388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1389 = {1{$random}};
  mem_1389 = _RAND_1389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1390 = {1{$random}};
  mem_1390 = _RAND_1390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1391 = {1{$random}};
  mem_1391 = _RAND_1391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1392 = {1{$random}};
  mem_1392 = _RAND_1392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1393 = {1{$random}};
  mem_1393 = _RAND_1393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1394 = {1{$random}};
  mem_1394 = _RAND_1394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1395 = {1{$random}};
  mem_1395 = _RAND_1395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1396 = {1{$random}};
  mem_1396 = _RAND_1396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1397 = {1{$random}};
  mem_1397 = _RAND_1397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1398 = {1{$random}};
  mem_1398 = _RAND_1398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1399 = {1{$random}};
  mem_1399 = _RAND_1399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1400 = {1{$random}};
  mem_1400 = _RAND_1400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1401 = {1{$random}};
  mem_1401 = _RAND_1401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1402 = {1{$random}};
  mem_1402 = _RAND_1402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1403 = {1{$random}};
  mem_1403 = _RAND_1403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1404 = {1{$random}};
  mem_1404 = _RAND_1404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1405 = {1{$random}};
  mem_1405 = _RAND_1405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1406 = {1{$random}};
  mem_1406 = _RAND_1406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1407 = {1{$random}};
  mem_1407 = _RAND_1407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1408 = {1{$random}};
  mem_1408 = _RAND_1408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1409 = {1{$random}};
  mem_1409 = _RAND_1409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1410 = {1{$random}};
  mem_1410 = _RAND_1410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1411 = {1{$random}};
  mem_1411 = _RAND_1411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1412 = {1{$random}};
  mem_1412 = _RAND_1412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1413 = {1{$random}};
  mem_1413 = _RAND_1413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1414 = {1{$random}};
  mem_1414 = _RAND_1414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1415 = {1{$random}};
  mem_1415 = _RAND_1415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1416 = {1{$random}};
  mem_1416 = _RAND_1416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1417 = {1{$random}};
  mem_1417 = _RAND_1417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1418 = {1{$random}};
  mem_1418 = _RAND_1418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1419 = {1{$random}};
  mem_1419 = _RAND_1419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1420 = {1{$random}};
  mem_1420 = _RAND_1420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1421 = {1{$random}};
  mem_1421 = _RAND_1421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1422 = {1{$random}};
  mem_1422 = _RAND_1422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1423 = {1{$random}};
  mem_1423 = _RAND_1423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1424 = {1{$random}};
  mem_1424 = _RAND_1424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1425 = {1{$random}};
  mem_1425 = _RAND_1425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1426 = {1{$random}};
  mem_1426 = _RAND_1426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1427 = {1{$random}};
  mem_1427 = _RAND_1427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1428 = {1{$random}};
  mem_1428 = _RAND_1428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1429 = {1{$random}};
  mem_1429 = _RAND_1429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1430 = {1{$random}};
  mem_1430 = _RAND_1430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1431 = {1{$random}};
  mem_1431 = _RAND_1431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1432 = {1{$random}};
  mem_1432 = _RAND_1432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1433 = {1{$random}};
  mem_1433 = _RAND_1433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1434 = {1{$random}};
  mem_1434 = _RAND_1434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1435 = {1{$random}};
  mem_1435 = _RAND_1435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1436 = {1{$random}};
  mem_1436 = _RAND_1436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1437 = {1{$random}};
  mem_1437 = _RAND_1437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1438 = {1{$random}};
  mem_1438 = _RAND_1438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1439 = {1{$random}};
  mem_1439 = _RAND_1439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1440 = {1{$random}};
  mem_1440 = _RAND_1440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1441 = {1{$random}};
  mem_1441 = _RAND_1441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1442 = {1{$random}};
  mem_1442 = _RAND_1442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1443 = {1{$random}};
  mem_1443 = _RAND_1443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1444 = {1{$random}};
  mem_1444 = _RAND_1444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1445 = {1{$random}};
  mem_1445 = _RAND_1445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1446 = {1{$random}};
  mem_1446 = _RAND_1446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1447 = {1{$random}};
  mem_1447 = _RAND_1447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1448 = {1{$random}};
  mem_1448 = _RAND_1448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1449 = {1{$random}};
  mem_1449 = _RAND_1449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1450 = {1{$random}};
  mem_1450 = _RAND_1450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1451 = {1{$random}};
  mem_1451 = _RAND_1451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1452 = {1{$random}};
  mem_1452 = _RAND_1452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1453 = {1{$random}};
  mem_1453 = _RAND_1453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1454 = {1{$random}};
  mem_1454 = _RAND_1454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1455 = {1{$random}};
  mem_1455 = _RAND_1455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1456 = {1{$random}};
  mem_1456 = _RAND_1456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1457 = {1{$random}};
  mem_1457 = _RAND_1457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1458 = {1{$random}};
  mem_1458 = _RAND_1458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1459 = {1{$random}};
  mem_1459 = _RAND_1459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1460 = {1{$random}};
  mem_1460 = _RAND_1460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1461 = {1{$random}};
  mem_1461 = _RAND_1461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1462 = {1{$random}};
  mem_1462 = _RAND_1462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1463 = {1{$random}};
  mem_1463 = _RAND_1463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1464 = {1{$random}};
  mem_1464 = _RAND_1464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1465 = {1{$random}};
  mem_1465 = _RAND_1465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1466 = {1{$random}};
  mem_1466 = _RAND_1466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1467 = {1{$random}};
  mem_1467 = _RAND_1467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1468 = {1{$random}};
  mem_1468 = _RAND_1468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1469 = {1{$random}};
  mem_1469 = _RAND_1469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1470 = {1{$random}};
  mem_1470 = _RAND_1470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1471 = {1{$random}};
  mem_1471 = _RAND_1471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1472 = {1{$random}};
  mem_1472 = _RAND_1472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1473 = {1{$random}};
  mem_1473 = _RAND_1473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1474 = {1{$random}};
  mem_1474 = _RAND_1474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1475 = {1{$random}};
  mem_1475 = _RAND_1475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1476 = {1{$random}};
  mem_1476 = _RAND_1476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1477 = {1{$random}};
  mem_1477 = _RAND_1477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1478 = {1{$random}};
  mem_1478 = _RAND_1478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1479 = {1{$random}};
  mem_1479 = _RAND_1479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1480 = {1{$random}};
  mem_1480 = _RAND_1480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1481 = {1{$random}};
  mem_1481 = _RAND_1481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1482 = {1{$random}};
  mem_1482 = _RAND_1482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1483 = {1{$random}};
  mem_1483 = _RAND_1483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1484 = {1{$random}};
  mem_1484 = _RAND_1484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1485 = {1{$random}};
  mem_1485 = _RAND_1485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1486 = {1{$random}};
  mem_1486 = _RAND_1486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1487 = {1{$random}};
  mem_1487 = _RAND_1487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1488 = {1{$random}};
  mem_1488 = _RAND_1488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1489 = {1{$random}};
  mem_1489 = _RAND_1489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1490 = {1{$random}};
  mem_1490 = _RAND_1490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1491 = {1{$random}};
  mem_1491 = _RAND_1491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1492 = {1{$random}};
  mem_1492 = _RAND_1492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1493 = {1{$random}};
  mem_1493 = _RAND_1493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1494 = {1{$random}};
  mem_1494 = _RAND_1494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1495 = {1{$random}};
  mem_1495 = _RAND_1495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1496 = {1{$random}};
  mem_1496 = _RAND_1496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1497 = {1{$random}};
  mem_1497 = _RAND_1497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1498 = {1{$random}};
  mem_1498 = _RAND_1498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1499 = {1{$random}};
  mem_1499 = _RAND_1499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1500 = {1{$random}};
  mem_1500 = _RAND_1500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1501 = {1{$random}};
  mem_1501 = _RAND_1501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1502 = {1{$random}};
  mem_1502 = _RAND_1502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1503 = {1{$random}};
  mem_1503 = _RAND_1503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1504 = {1{$random}};
  mem_1504 = _RAND_1504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1505 = {1{$random}};
  mem_1505 = _RAND_1505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1506 = {1{$random}};
  mem_1506 = _RAND_1506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1507 = {1{$random}};
  mem_1507 = _RAND_1507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1508 = {1{$random}};
  mem_1508 = _RAND_1508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1509 = {1{$random}};
  mem_1509 = _RAND_1509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1510 = {1{$random}};
  mem_1510 = _RAND_1510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1511 = {1{$random}};
  mem_1511 = _RAND_1511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1512 = {1{$random}};
  mem_1512 = _RAND_1512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1513 = {1{$random}};
  mem_1513 = _RAND_1513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1514 = {1{$random}};
  mem_1514 = _RAND_1514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1515 = {1{$random}};
  mem_1515 = _RAND_1515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1516 = {1{$random}};
  mem_1516 = _RAND_1516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1517 = {1{$random}};
  mem_1517 = _RAND_1517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1518 = {1{$random}};
  mem_1518 = _RAND_1518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1519 = {1{$random}};
  mem_1519 = _RAND_1519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1520 = {1{$random}};
  mem_1520 = _RAND_1520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1521 = {1{$random}};
  mem_1521 = _RAND_1521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1522 = {1{$random}};
  mem_1522 = _RAND_1522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1523 = {1{$random}};
  mem_1523 = _RAND_1523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1524 = {1{$random}};
  mem_1524 = _RAND_1524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1525 = {1{$random}};
  mem_1525 = _RAND_1525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1526 = {1{$random}};
  mem_1526 = _RAND_1526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1527 = {1{$random}};
  mem_1527 = _RAND_1527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1528 = {1{$random}};
  mem_1528 = _RAND_1528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1529 = {1{$random}};
  mem_1529 = _RAND_1529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1530 = {1{$random}};
  mem_1530 = _RAND_1530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1531 = {1{$random}};
  mem_1531 = _RAND_1531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1532 = {1{$random}};
  mem_1532 = _RAND_1532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1533 = {1{$random}};
  mem_1533 = _RAND_1533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1534 = {1{$random}};
  mem_1534 = _RAND_1534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1535 = {1{$random}};
  mem_1535 = _RAND_1535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1536 = {1{$random}};
  mem_1536 = _RAND_1536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1537 = {1{$random}};
  mem_1537 = _RAND_1537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1538 = {1{$random}};
  mem_1538 = _RAND_1538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1539 = {1{$random}};
  mem_1539 = _RAND_1539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1540 = {1{$random}};
  mem_1540 = _RAND_1540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1541 = {1{$random}};
  mem_1541 = _RAND_1541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1542 = {1{$random}};
  mem_1542 = _RAND_1542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1543 = {1{$random}};
  mem_1543 = _RAND_1543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1544 = {1{$random}};
  mem_1544 = _RAND_1544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1545 = {1{$random}};
  mem_1545 = _RAND_1545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1546 = {1{$random}};
  mem_1546 = _RAND_1546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1547 = {1{$random}};
  mem_1547 = _RAND_1547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1548 = {1{$random}};
  mem_1548 = _RAND_1548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1549 = {1{$random}};
  mem_1549 = _RAND_1549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1550 = {1{$random}};
  mem_1550 = _RAND_1550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1551 = {1{$random}};
  mem_1551 = _RAND_1551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1552 = {1{$random}};
  mem_1552 = _RAND_1552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1553 = {1{$random}};
  mem_1553 = _RAND_1553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1554 = {1{$random}};
  mem_1554 = _RAND_1554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1555 = {1{$random}};
  mem_1555 = _RAND_1555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1556 = {1{$random}};
  mem_1556 = _RAND_1556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1557 = {1{$random}};
  mem_1557 = _RAND_1557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1558 = {1{$random}};
  mem_1558 = _RAND_1558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1559 = {1{$random}};
  mem_1559 = _RAND_1559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1560 = {1{$random}};
  mem_1560 = _RAND_1560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1561 = {1{$random}};
  mem_1561 = _RAND_1561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1562 = {1{$random}};
  mem_1562 = _RAND_1562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1563 = {1{$random}};
  mem_1563 = _RAND_1563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1564 = {1{$random}};
  mem_1564 = _RAND_1564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1565 = {1{$random}};
  mem_1565 = _RAND_1565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1566 = {1{$random}};
  mem_1566 = _RAND_1566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1567 = {1{$random}};
  mem_1567 = _RAND_1567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1568 = {1{$random}};
  mem_1568 = _RAND_1568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1569 = {1{$random}};
  mem_1569 = _RAND_1569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1570 = {1{$random}};
  mem_1570 = _RAND_1570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1571 = {1{$random}};
  mem_1571 = _RAND_1571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1572 = {1{$random}};
  mem_1572 = _RAND_1572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1573 = {1{$random}};
  mem_1573 = _RAND_1573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1574 = {1{$random}};
  mem_1574 = _RAND_1574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1575 = {1{$random}};
  mem_1575 = _RAND_1575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1576 = {1{$random}};
  mem_1576 = _RAND_1576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1577 = {1{$random}};
  mem_1577 = _RAND_1577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1578 = {1{$random}};
  mem_1578 = _RAND_1578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1579 = {1{$random}};
  mem_1579 = _RAND_1579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1580 = {1{$random}};
  mem_1580 = _RAND_1580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1581 = {1{$random}};
  mem_1581 = _RAND_1581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1582 = {1{$random}};
  mem_1582 = _RAND_1582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1583 = {1{$random}};
  mem_1583 = _RAND_1583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1584 = {1{$random}};
  mem_1584 = _RAND_1584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1585 = {1{$random}};
  mem_1585 = _RAND_1585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1586 = {1{$random}};
  mem_1586 = _RAND_1586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1587 = {1{$random}};
  mem_1587 = _RAND_1587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1588 = {1{$random}};
  mem_1588 = _RAND_1588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1589 = {1{$random}};
  mem_1589 = _RAND_1589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1590 = {1{$random}};
  mem_1590 = _RAND_1590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1591 = {1{$random}};
  mem_1591 = _RAND_1591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1592 = {1{$random}};
  mem_1592 = _RAND_1592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1593 = {1{$random}};
  mem_1593 = _RAND_1593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1594 = {1{$random}};
  mem_1594 = _RAND_1594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1595 = {1{$random}};
  mem_1595 = _RAND_1595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1596 = {1{$random}};
  mem_1596 = _RAND_1596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1597 = {1{$random}};
  mem_1597 = _RAND_1597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1598 = {1{$random}};
  mem_1598 = _RAND_1598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1599 = {1{$random}};
  mem_1599 = _RAND_1599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1600 = {1{$random}};
  mem_1600 = _RAND_1600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1601 = {1{$random}};
  mem_1601 = _RAND_1601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1602 = {1{$random}};
  mem_1602 = _RAND_1602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1603 = {1{$random}};
  mem_1603 = _RAND_1603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1604 = {1{$random}};
  mem_1604 = _RAND_1604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1605 = {1{$random}};
  mem_1605 = _RAND_1605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1606 = {1{$random}};
  mem_1606 = _RAND_1606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1607 = {1{$random}};
  mem_1607 = _RAND_1607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1608 = {1{$random}};
  mem_1608 = _RAND_1608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1609 = {1{$random}};
  mem_1609 = _RAND_1609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1610 = {1{$random}};
  mem_1610 = _RAND_1610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1611 = {1{$random}};
  mem_1611 = _RAND_1611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1612 = {1{$random}};
  mem_1612 = _RAND_1612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1613 = {1{$random}};
  mem_1613 = _RAND_1613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1614 = {1{$random}};
  mem_1614 = _RAND_1614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1615 = {1{$random}};
  mem_1615 = _RAND_1615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1616 = {1{$random}};
  mem_1616 = _RAND_1616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1617 = {1{$random}};
  mem_1617 = _RAND_1617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1618 = {1{$random}};
  mem_1618 = _RAND_1618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1619 = {1{$random}};
  mem_1619 = _RAND_1619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1620 = {1{$random}};
  mem_1620 = _RAND_1620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1621 = {1{$random}};
  mem_1621 = _RAND_1621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1622 = {1{$random}};
  mem_1622 = _RAND_1622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1623 = {1{$random}};
  mem_1623 = _RAND_1623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1624 = {1{$random}};
  mem_1624 = _RAND_1624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1625 = {1{$random}};
  mem_1625 = _RAND_1625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1626 = {1{$random}};
  mem_1626 = _RAND_1626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1627 = {1{$random}};
  mem_1627 = _RAND_1627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1628 = {1{$random}};
  mem_1628 = _RAND_1628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1629 = {1{$random}};
  mem_1629 = _RAND_1629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1630 = {1{$random}};
  mem_1630 = _RAND_1630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1631 = {1{$random}};
  mem_1631 = _RAND_1631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1632 = {1{$random}};
  mem_1632 = _RAND_1632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1633 = {1{$random}};
  mem_1633 = _RAND_1633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1634 = {1{$random}};
  mem_1634 = _RAND_1634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1635 = {1{$random}};
  mem_1635 = _RAND_1635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1636 = {1{$random}};
  mem_1636 = _RAND_1636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1637 = {1{$random}};
  mem_1637 = _RAND_1637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1638 = {1{$random}};
  mem_1638 = _RAND_1638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1639 = {1{$random}};
  mem_1639 = _RAND_1639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1640 = {1{$random}};
  mem_1640 = _RAND_1640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1641 = {1{$random}};
  mem_1641 = _RAND_1641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1642 = {1{$random}};
  mem_1642 = _RAND_1642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1643 = {1{$random}};
  mem_1643 = _RAND_1643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1644 = {1{$random}};
  mem_1644 = _RAND_1644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1645 = {1{$random}};
  mem_1645 = _RAND_1645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1646 = {1{$random}};
  mem_1646 = _RAND_1646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1647 = {1{$random}};
  mem_1647 = _RAND_1647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1648 = {1{$random}};
  mem_1648 = _RAND_1648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1649 = {1{$random}};
  mem_1649 = _RAND_1649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1650 = {1{$random}};
  mem_1650 = _RAND_1650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1651 = {1{$random}};
  mem_1651 = _RAND_1651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1652 = {1{$random}};
  mem_1652 = _RAND_1652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1653 = {1{$random}};
  mem_1653 = _RAND_1653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1654 = {1{$random}};
  mem_1654 = _RAND_1654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1655 = {1{$random}};
  mem_1655 = _RAND_1655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1656 = {1{$random}};
  mem_1656 = _RAND_1656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1657 = {1{$random}};
  mem_1657 = _RAND_1657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1658 = {1{$random}};
  mem_1658 = _RAND_1658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1659 = {1{$random}};
  mem_1659 = _RAND_1659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1660 = {1{$random}};
  mem_1660 = _RAND_1660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1661 = {1{$random}};
  mem_1661 = _RAND_1661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1662 = {1{$random}};
  mem_1662 = _RAND_1662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1663 = {1{$random}};
  mem_1663 = _RAND_1663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1664 = {1{$random}};
  mem_1664 = _RAND_1664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1665 = {1{$random}};
  mem_1665 = _RAND_1665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1666 = {1{$random}};
  mem_1666 = _RAND_1666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1667 = {1{$random}};
  mem_1667 = _RAND_1667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1668 = {1{$random}};
  mem_1668 = _RAND_1668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1669 = {1{$random}};
  mem_1669 = _RAND_1669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1670 = {1{$random}};
  mem_1670 = _RAND_1670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1671 = {1{$random}};
  mem_1671 = _RAND_1671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1672 = {1{$random}};
  mem_1672 = _RAND_1672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1673 = {1{$random}};
  mem_1673 = _RAND_1673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1674 = {1{$random}};
  mem_1674 = _RAND_1674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1675 = {1{$random}};
  mem_1675 = _RAND_1675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1676 = {1{$random}};
  mem_1676 = _RAND_1676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1677 = {1{$random}};
  mem_1677 = _RAND_1677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1678 = {1{$random}};
  mem_1678 = _RAND_1678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1679 = {1{$random}};
  mem_1679 = _RAND_1679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1680 = {1{$random}};
  mem_1680 = _RAND_1680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1681 = {1{$random}};
  mem_1681 = _RAND_1681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1682 = {1{$random}};
  mem_1682 = _RAND_1682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1683 = {1{$random}};
  mem_1683 = _RAND_1683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1684 = {1{$random}};
  mem_1684 = _RAND_1684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1685 = {1{$random}};
  mem_1685 = _RAND_1685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1686 = {1{$random}};
  mem_1686 = _RAND_1686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1687 = {1{$random}};
  mem_1687 = _RAND_1687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1688 = {1{$random}};
  mem_1688 = _RAND_1688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1689 = {1{$random}};
  mem_1689 = _RAND_1689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1690 = {1{$random}};
  mem_1690 = _RAND_1690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1691 = {1{$random}};
  mem_1691 = _RAND_1691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1692 = {1{$random}};
  mem_1692 = _RAND_1692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1693 = {1{$random}};
  mem_1693 = _RAND_1693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1694 = {1{$random}};
  mem_1694 = _RAND_1694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1695 = {1{$random}};
  mem_1695 = _RAND_1695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1696 = {1{$random}};
  mem_1696 = _RAND_1696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1697 = {1{$random}};
  mem_1697 = _RAND_1697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1698 = {1{$random}};
  mem_1698 = _RAND_1698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1699 = {1{$random}};
  mem_1699 = _RAND_1699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1700 = {1{$random}};
  mem_1700 = _RAND_1700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1701 = {1{$random}};
  mem_1701 = _RAND_1701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1702 = {1{$random}};
  mem_1702 = _RAND_1702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1703 = {1{$random}};
  mem_1703 = _RAND_1703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1704 = {1{$random}};
  mem_1704 = _RAND_1704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1705 = {1{$random}};
  mem_1705 = _RAND_1705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1706 = {1{$random}};
  mem_1706 = _RAND_1706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1707 = {1{$random}};
  mem_1707 = _RAND_1707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1708 = {1{$random}};
  mem_1708 = _RAND_1708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1709 = {1{$random}};
  mem_1709 = _RAND_1709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1710 = {1{$random}};
  mem_1710 = _RAND_1710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1711 = {1{$random}};
  mem_1711 = _RAND_1711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1712 = {1{$random}};
  mem_1712 = _RAND_1712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1713 = {1{$random}};
  mem_1713 = _RAND_1713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1714 = {1{$random}};
  mem_1714 = _RAND_1714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1715 = {1{$random}};
  mem_1715 = _RAND_1715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1716 = {1{$random}};
  mem_1716 = _RAND_1716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1717 = {1{$random}};
  mem_1717 = _RAND_1717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1718 = {1{$random}};
  mem_1718 = _RAND_1718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1719 = {1{$random}};
  mem_1719 = _RAND_1719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1720 = {1{$random}};
  mem_1720 = _RAND_1720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1721 = {1{$random}};
  mem_1721 = _RAND_1721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1722 = {1{$random}};
  mem_1722 = _RAND_1722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1723 = {1{$random}};
  mem_1723 = _RAND_1723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1724 = {1{$random}};
  mem_1724 = _RAND_1724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1725 = {1{$random}};
  mem_1725 = _RAND_1725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1726 = {1{$random}};
  mem_1726 = _RAND_1726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1727 = {1{$random}};
  mem_1727 = _RAND_1727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1728 = {1{$random}};
  mem_1728 = _RAND_1728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1729 = {1{$random}};
  mem_1729 = _RAND_1729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1730 = {1{$random}};
  mem_1730 = _RAND_1730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1731 = {1{$random}};
  mem_1731 = _RAND_1731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1732 = {1{$random}};
  mem_1732 = _RAND_1732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1733 = {1{$random}};
  mem_1733 = _RAND_1733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1734 = {1{$random}};
  mem_1734 = _RAND_1734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1735 = {1{$random}};
  mem_1735 = _RAND_1735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1736 = {1{$random}};
  mem_1736 = _RAND_1736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1737 = {1{$random}};
  mem_1737 = _RAND_1737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1738 = {1{$random}};
  mem_1738 = _RAND_1738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1739 = {1{$random}};
  mem_1739 = _RAND_1739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1740 = {1{$random}};
  mem_1740 = _RAND_1740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1741 = {1{$random}};
  mem_1741 = _RAND_1741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1742 = {1{$random}};
  mem_1742 = _RAND_1742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1743 = {1{$random}};
  mem_1743 = _RAND_1743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1744 = {1{$random}};
  mem_1744 = _RAND_1744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1745 = {1{$random}};
  mem_1745 = _RAND_1745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1746 = {1{$random}};
  mem_1746 = _RAND_1746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1747 = {1{$random}};
  mem_1747 = _RAND_1747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1748 = {1{$random}};
  mem_1748 = _RAND_1748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1749 = {1{$random}};
  mem_1749 = _RAND_1749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1750 = {1{$random}};
  mem_1750 = _RAND_1750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1751 = {1{$random}};
  mem_1751 = _RAND_1751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1752 = {1{$random}};
  mem_1752 = _RAND_1752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1753 = {1{$random}};
  mem_1753 = _RAND_1753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1754 = {1{$random}};
  mem_1754 = _RAND_1754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1755 = {1{$random}};
  mem_1755 = _RAND_1755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1756 = {1{$random}};
  mem_1756 = _RAND_1756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1757 = {1{$random}};
  mem_1757 = _RAND_1757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1758 = {1{$random}};
  mem_1758 = _RAND_1758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1759 = {1{$random}};
  mem_1759 = _RAND_1759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1760 = {1{$random}};
  mem_1760 = _RAND_1760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1761 = {1{$random}};
  mem_1761 = _RAND_1761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1762 = {1{$random}};
  mem_1762 = _RAND_1762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1763 = {1{$random}};
  mem_1763 = _RAND_1763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1764 = {1{$random}};
  mem_1764 = _RAND_1764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1765 = {1{$random}};
  mem_1765 = _RAND_1765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1766 = {1{$random}};
  mem_1766 = _RAND_1766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1767 = {1{$random}};
  mem_1767 = _RAND_1767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1768 = {1{$random}};
  mem_1768 = _RAND_1768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1769 = {1{$random}};
  mem_1769 = _RAND_1769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1770 = {1{$random}};
  mem_1770 = _RAND_1770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1771 = {1{$random}};
  mem_1771 = _RAND_1771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1772 = {1{$random}};
  mem_1772 = _RAND_1772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1773 = {1{$random}};
  mem_1773 = _RAND_1773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1774 = {1{$random}};
  mem_1774 = _RAND_1774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1775 = {1{$random}};
  mem_1775 = _RAND_1775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1776 = {1{$random}};
  mem_1776 = _RAND_1776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1777 = {1{$random}};
  mem_1777 = _RAND_1777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1778 = {1{$random}};
  mem_1778 = _RAND_1778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1779 = {1{$random}};
  mem_1779 = _RAND_1779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1780 = {1{$random}};
  mem_1780 = _RAND_1780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1781 = {1{$random}};
  mem_1781 = _RAND_1781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1782 = {1{$random}};
  mem_1782 = _RAND_1782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1783 = {1{$random}};
  mem_1783 = _RAND_1783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1784 = {1{$random}};
  mem_1784 = _RAND_1784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1785 = {1{$random}};
  mem_1785 = _RAND_1785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1786 = {1{$random}};
  mem_1786 = _RAND_1786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1787 = {1{$random}};
  mem_1787 = _RAND_1787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1788 = {1{$random}};
  mem_1788 = _RAND_1788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1789 = {1{$random}};
  mem_1789 = _RAND_1789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1790 = {1{$random}};
  mem_1790 = _RAND_1790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1791 = {1{$random}};
  mem_1791 = _RAND_1791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1792 = {1{$random}};
  mem_1792 = _RAND_1792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1793 = {1{$random}};
  mem_1793 = _RAND_1793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1794 = {1{$random}};
  mem_1794 = _RAND_1794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1795 = {1{$random}};
  mem_1795 = _RAND_1795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1796 = {1{$random}};
  mem_1796 = _RAND_1796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1797 = {1{$random}};
  mem_1797 = _RAND_1797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1798 = {1{$random}};
  mem_1798 = _RAND_1798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1799 = {1{$random}};
  mem_1799 = _RAND_1799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1800 = {1{$random}};
  mem_1800 = _RAND_1800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1801 = {1{$random}};
  mem_1801 = _RAND_1801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1802 = {1{$random}};
  mem_1802 = _RAND_1802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1803 = {1{$random}};
  mem_1803 = _RAND_1803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1804 = {1{$random}};
  mem_1804 = _RAND_1804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1805 = {1{$random}};
  mem_1805 = _RAND_1805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1806 = {1{$random}};
  mem_1806 = _RAND_1806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1807 = {1{$random}};
  mem_1807 = _RAND_1807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1808 = {1{$random}};
  mem_1808 = _RAND_1808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1809 = {1{$random}};
  mem_1809 = _RAND_1809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1810 = {1{$random}};
  mem_1810 = _RAND_1810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1811 = {1{$random}};
  mem_1811 = _RAND_1811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1812 = {1{$random}};
  mem_1812 = _RAND_1812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1813 = {1{$random}};
  mem_1813 = _RAND_1813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1814 = {1{$random}};
  mem_1814 = _RAND_1814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1815 = {1{$random}};
  mem_1815 = _RAND_1815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1816 = {1{$random}};
  mem_1816 = _RAND_1816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1817 = {1{$random}};
  mem_1817 = _RAND_1817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1818 = {1{$random}};
  mem_1818 = _RAND_1818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1819 = {1{$random}};
  mem_1819 = _RAND_1819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1820 = {1{$random}};
  mem_1820 = _RAND_1820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1821 = {1{$random}};
  mem_1821 = _RAND_1821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1822 = {1{$random}};
  mem_1822 = _RAND_1822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1823 = {1{$random}};
  mem_1823 = _RAND_1823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1824 = {1{$random}};
  mem_1824 = _RAND_1824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1825 = {1{$random}};
  mem_1825 = _RAND_1825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1826 = {1{$random}};
  mem_1826 = _RAND_1826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1827 = {1{$random}};
  mem_1827 = _RAND_1827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1828 = {1{$random}};
  mem_1828 = _RAND_1828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1829 = {1{$random}};
  mem_1829 = _RAND_1829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1830 = {1{$random}};
  mem_1830 = _RAND_1830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1831 = {1{$random}};
  mem_1831 = _RAND_1831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1832 = {1{$random}};
  mem_1832 = _RAND_1832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1833 = {1{$random}};
  mem_1833 = _RAND_1833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1834 = {1{$random}};
  mem_1834 = _RAND_1834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1835 = {1{$random}};
  mem_1835 = _RAND_1835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1836 = {1{$random}};
  mem_1836 = _RAND_1836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1837 = {1{$random}};
  mem_1837 = _RAND_1837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1838 = {1{$random}};
  mem_1838 = _RAND_1838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1839 = {1{$random}};
  mem_1839 = _RAND_1839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1840 = {1{$random}};
  mem_1840 = _RAND_1840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1841 = {1{$random}};
  mem_1841 = _RAND_1841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1842 = {1{$random}};
  mem_1842 = _RAND_1842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1843 = {1{$random}};
  mem_1843 = _RAND_1843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1844 = {1{$random}};
  mem_1844 = _RAND_1844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1845 = {1{$random}};
  mem_1845 = _RAND_1845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1846 = {1{$random}};
  mem_1846 = _RAND_1846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1847 = {1{$random}};
  mem_1847 = _RAND_1847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1848 = {1{$random}};
  mem_1848 = _RAND_1848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1849 = {1{$random}};
  mem_1849 = _RAND_1849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1850 = {1{$random}};
  mem_1850 = _RAND_1850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1851 = {1{$random}};
  mem_1851 = _RAND_1851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1852 = {1{$random}};
  mem_1852 = _RAND_1852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1853 = {1{$random}};
  mem_1853 = _RAND_1853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1854 = {1{$random}};
  mem_1854 = _RAND_1854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1855 = {1{$random}};
  mem_1855 = _RAND_1855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1856 = {1{$random}};
  mem_1856 = _RAND_1856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1857 = {1{$random}};
  mem_1857 = _RAND_1857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1858 = {1{$random}};
  mem_1858 = _RAND_1858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1859 = {1{$random}};
  mem_1859 = _RAND_1859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1860 = {1{$random}};
  mem_1860 = _RAND_1860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1861 = {1{$random}};
  mem_1861 = _RAND_1861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1862 = {1{$random}};
  mem_1862 = _RAND_1862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1863 = {1{$random}};
  mem_1863 = _RAND_1863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1864 = {1{$random}};
  mem_1864 = _RAND_1864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1865 = {1{$random}};
  mem_1865 = _RAND_1865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1866 = {1{$random}};
  mem_1866 = _RAND_1866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1867 = {1{$random}};
  mem_1867 = _RAND_1867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1868 = {1{$random}};
  mem_1868 = _RAND_1868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1869 = {1{$random}};
  mem_1869 = _RAND_1869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1870 = {1{$random}};
  mem_1870 = _RAND_1870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1871 = {1{$random}};
  mem_1871 = _RAND_1871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1872 = {1{$random}};
  mem_1872 = _RAND_1872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1873 = {1{$random}};
  mem_1873 = _RAND_1873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1874 = {1{$random}};
  mem_1874 = _RAND_1874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1875 = {1{$random}};
  mem_1875 = _RAND_1875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1876 = {1{$random}};
  mem_1876 = _RAND_1876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1877 = {1{$random}};
  mem_1877 = _RAND_1877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1878 = {1{$random}};
  mem_1878 = _RAND_1878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1879 = {1{$random}};
  mem_1879 = _RAND_1879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1880 = {1{$random}};
  mem_1880 = _RAND_1880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1881 = {1{$random}};
  mem_1881 = _RAND_1881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1882 = {1{$random}};
  mem_1882 = _RAND_1882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1883 = {1{$random}};
  mem_1883 = _RAND_1883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1884 = {1{$random}};
  mem_1884 = _RAND_1884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1885 = {1{$random}};
  mem_1885 = _RAND_1885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1886 = {1{$random}};
  mem_1886 = _RAND_1886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1887 = {1{$random}};
  mem_1887 = _RAND_1887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1888 = {1{$random}};
  mem_1888 = _RAND_1888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1889 = {1{$random}};
  mem_1889 = _RAND_1889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1890 = {1{$random}};
  mem_1890 = _RAND_1890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1891 = {1{$random}};
  mem_1891 = _RAND_1891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1892 = {1{$random}};
  mem_1892 = _RAND_1892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1893 = {1{$random}};
  mem_1893 = _RAND_1893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1894 = {1{$random}};
  mem_1894 = _RAND_1894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1895 = {1{$random}};
  mem_1895 = _RAND_1895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1896 = {1{$random}};
  mem_1896 = _RAND_1896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1897 = {1{$random}};
  mem_1897 = _RAND_1897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1898 = {1{$random}};
  mem_1898 = _RAND_1898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1899 = {1{$random}};
  mem_1899 = _RAND_1899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1900 = {1{$random}};
  mem_1900 = _RAND_1900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1901 = {1{$random}};
  mem_1901 = _RAND_1901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1902 = {1{$random}};
  mem_1902 = _RAND_1902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1903 = {1{$random}};
  mem_1903 = _RAND_1903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1904 = {1{$random}};
  mem_1904 = _RAND_1904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1905 = {1{$random}};
  mem_1905 = _RAND_1905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1906 = {1{$random}};
  mem_1906 = _RAND_1906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1907 = {1{$random}};
  mem_1907 = _RAND_1907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1908 = {1{$random}};
  mem_1908 = _RAND_1908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1909 = {1{$random}};
  mem_1909 = _RAND_1909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1910 = {1{$random}};
  mem_1910 = _RAND_1910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1911 = {1{$random}};
  mem_1911 = _RAND_1911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1912 = {1{$random}};
  mem_1912 = _RAND_1912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1913 = {1{$random}};
  mem_1913 = _RAND_1913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1914 = {1{$random}};
  mem_1914 = _RAND_1914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1915 = {1{$random}};
  mem_1915 = _RAND_1915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1916 = {1{$random}};
  mem_1916 = _RAND_1916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1917 = {1{$random}};
  mem_1917 = _RAND_1917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1918 = {1{$random}};
  mem_1918 = _RAND_1918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1919 = {1{$random}};
  mem_1919 = _RAND_1919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1920 = {1{$random}};
  mem_1920 = _RAND_1920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1921 = {1{$random}};
  mem_1921 = _RAND_1921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1922 = {1{$random}};
  mem_1922 = _RAND_1922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1923 = {1{$random}};
  mem_1923 = _RAND_1923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1924 = {1{$random}};
  mem_1924 = _RAND_1924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1925 = {1{$random}};
  mem_1925 = _RAND_1925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1926 = {1{$random}};
  mem_1926 = _RAND_1926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1927 = {1{$random}};
  mem_1927 = _RAND_1927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1928 = {1{$random}};
  mem_1928 = _RAND_1928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1929 = {1{$random}};
  mem_1929 = _RAND_1929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1930 = {1{$random}};
  mem_1930 = _RAND_1930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1931 = {1{$random}};
  mem_1931 = _RAND_1931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1932 = {1{$random}};
  mem_1932 = _RAND_1932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1933 = {1{$random}};
  mem_1933 = _RAND_1933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1934 = {1{$random}};
  mem_1934 = _RAND_1934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1935 = {1{$random}};
  mem_1935 = _RAND_1935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1936 = {1{$random}};
  mem_1936 = _RAND_1936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1937 = {1{$random}};
  mem_1937 = _RAND_1937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1938 = {1{$random}};
  mem_1938 = _RAND_1938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1939 = {1{$random}};
  mem_1939 = _RAND_1939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1940 = {1{$random}};
  mem_1940 = _RAND_1940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1941 = {1{$random}};
  mem_1941 = _RAND_1941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1942 = {1{$random}};
  mem_1942 = _RAND_1942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1943 = {1{$random}};
  mem_1943 = _RAND_1943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1944 = {1{$random}};
  mem_1944 = _RAND_1944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1945 = {1{$random}};
  mem_1945 = _RAND_1945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1946 = {1{$random}};
  mem_1946 = _RAND_1946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1947 = {1{$random}};
  mem_1947 = _RAND_1947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1948 = {1{$random}};
  mem_1948 = _RAND_1948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1949 = {1{$random}};
  mem_1949 = _RAND_1949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1950 = {1{$random}};
  mem_1950 = _RAND_1950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1951 = {1{$random}};
  mem_1951 = _RAND_1951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1952 = {1{$random}};
  mem_1952 = _RAND_1952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1953 = {1{$random}};
  mem_1953 = _RAND_1953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1954 = {1{$random}};
  mem_1954 = _RAND_1954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1955 = {1{$random}};
  mem_1955 = _RAND_1955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1956 = {1{$random}};
  mem_1956 = _RAND_1956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1957 = {1{$random}};
  mem_1957 = _RAND_1957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1958 = {1{$random}};
  mem_1958 = _RAND_1958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1959 = {1{$random}};
  mem_1959 = _RAND_1959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1960 = {1{$random}};
  mem_1960 = _RAND_1960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1961 = {1{$random}};
  mem_1961 = _RAND_1961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1962 = {1{$random}};
  mem_1962 = _RAND_1962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1963 = {1{$random}};
  mem_1963 = _RAND_1963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1964 = {1{$random}};
  mem_1964 = _RAND_1964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1965 = {1{$random}};
  mem_1965 = _RAND_1965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1966 = {1{$random}};
  mem_1966 = _RAND_1966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1967 = {1{$random}};
  mem_1967 = _RAND_1967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1968 = {1{$random}};
  mem_1968 = _RAND_1968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1969 = {1{$random}};
  mem_1969 = _RAND_1969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1970 = {1{$random}};
  mem_1970 = _RAND_1970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1971 = {1{$random}};
  mem_1971 = _RAND_1971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1972 = {1{$random}};
  mem_1972 = _RAND_1972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1973 = {1{$random}};
  mem_1973 = _RAND_1973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1974 = {1{$random}};
  mem_1974 = _RAND_1974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1975 = {1{$random}};
  mem_1975 = _RAND_1975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1976 = {1{$random}};
  mem_1976 = _RAND_1976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1977 = {1{$random}};
  mem_1977 = _RAND_1977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1978 = {1{$random}};
  mem_1978 = _RAND_1978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1979 = {1{$random}};
  mem_1979 = _RAND_1979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1980 = {1{$random}};
  mem_1980 = _RAND_1980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1981 = {1{$random}};
  mem_1981 = _RAND_1981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1982 = {1{$random}};
  mem_1982 = _RAND_1982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1983 = {1{$random}};
  mem_1983 = _RAND_1983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1984 = {1{$random}};
  mem_1984 = _RAND_1984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1985 = {1{$random}};
  mem_1985 = _RAND_1985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1986 = {1{$random}};
  mem_1986 = _RAND_1986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1987 = {1{$random}};
  mem_1987 = _RAND_1987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1988 = {1{$random}};
  mem_1988 = _RAND_1988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1989 = {1{$random}};
  mem_1989 = _RAND_1989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1990 = {1{$random}};
  mem_1990 = _RAND_1990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1991 = {1{$random}};
  mem_1991 = _RAND_1991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1992 = {1{$random}};
  mem_1992 = _RAND_1992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1993 = {1{$random}};
  mem_1993 = _RAND_1993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1994 = {1{$random}};
  mem_1994 = _RAND_1994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1995 = {1{$random}};
  mem_1995 = _RAND_1995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1996 = {1{$random}};
  mem_1996 = _RAND_1996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1997 = {1{$random}};
  mem_1997 = _RAND_1997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1998 = {1{$random}};
  mem_1998 = _RAND_1998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1999 = {1{$random}};
  mem_1999 = _RAND_1999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2000 = {1{$random}};
  mem_2000 = _RAND_2000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2001 = {1{$random}};
  mem_2001 = _RAND_2001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2002 = {1{$random}};
  mem_2002 = _RAND_2002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2003 = {1{$random}};
  mem_2003 = _RAND_2003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2004 = {1{$random}};
  mem_2004 = _RAND_2004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2005 = {1{$random}};
  mem_2005 = _RAND_2005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2006 = {1{$random}};
  mem_2006 = _RAND_2006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2007 = {1{$random}};
  mem_2007 = _RAND_2007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2008 = {1{$random}};
  mem_2008 = _RAND_2008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2009 = {1{$random}};
  mem_2009 = _RAND_2009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2010 = {1{$random}};
  mem_2010 = _RAND_2010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2011 = {1{$random}};
  mem_2011 = _RAND_2011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2012 = {1{$random}};
  mem_2012 = _RAND_2012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2013 = {1{$random}};
  mem_2013 = _RAND_2013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2014 = {1{$random}};
  mem_2014 = _RAND_2014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2015 = {1{$random}};
  mem_2015 = _RAND_2015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2016 = {1{$random}};
  mem_2016 = _RAND_2016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2017 = {1{$random}};
  mem_2017 = _RAND_2017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2018 = {1{$random}};
  mem_2018 = _RAND_2018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2019 = {1{$random}};
  mem_2019 = _RAND_2019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2020 = {1{$random}};
  mem_2020 = _RAND_2020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2021 = {1{$random}};
  mem_2021 = _RAND_2021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2022 = {1{$random}};
  mem_2022 = _RAND_2022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2023 = {1{$random}};
  mem_2023 = _RAND_2023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2024 = {1{$random}};
  mem_2024 = _RAND_2024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2025 = {1{$random}};
  mem_2025 = _RAND_2025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2026 = {1{$random}};
  mem_2026 = _RAND_2026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2027 = {1{$random}};
  mem_2027 = _RAND_2027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2028 = {1{$random}};
  mem_2028 = _RAND_2028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2029 = {1{$random}};
  mem_2029 = _RAND_2029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2030 = {1{$random}};
  mem_2030 = _RAND_2030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2031 = {1{$random}};
  mem_2031 = _RAND_2031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2032 = {1{$random}};
  mem_2032 = _RAND_2032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2033 = {1{$random}};
  mem_2033 = _RAND_2033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2034 = {1{$random}};
  mem_2034 = _RAND_2034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2035 = {1{$random}};
  mem_2035 = _RAND_2035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2036 = {1{$random}};
  mem_2036 = _RAND_2036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2037 = {1{$random}};
  mem_2037 = _RAND_2037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2038 = {1{$random}};
  mem_2038 = _RAND_2038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2039 = {1{$random}};
  mem_2039 = _RAND_2039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2040 = {1{$random}};
  mem_2040 = _RAND_2040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2041 = {1{$random}};
  mem_2041 = _RAND_2041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2042 = {1{$random}};
  mem_2042 = _RAND_2042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2043 = {1{$random}};
  mem_2043 = _RAND_2043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2044 = {1{$random}};
  mem_2044 = _RAND_2044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2045 = {1{$random}};
  mem_2045 = _RAND_2045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2046 = {1{$random}};
  mem_2046 = _RAND_2046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2047 = {1{$random}};
  mem_2047 = _RAND_2047[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      mem_0 <= 32'h2000537;
    end else begin
      if (11'h0 == _T_12323) begin
        mem_0 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1 <= 32'h450513;
    end else begin
      if (11'h1 == _T_12323) begin
        mem_1 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2 <= 32'h10f00593;
    end else begin
      if (11'h2 == _T_12323) begin
        mem_2 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_3 <= 32'hb52023;
    end else begin
      if (11'h3 == _T_12323) begin
        mem_3 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_4 <= 32'h450513;
    end else begin
      if (11'h4 == _T_12323) begin
        mem_4 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_5 <= 32'h4200593;
    end else begin
      if (11'h5 == _T_12323) begin
        mem_5 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_6 <= 32'hb52023;
    end else begin
      if (11'h6 == _T_12323) begin
        mem_6 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_7 <= 32'h6f00593;
    end else begin
      if (11'h7 == _T_12323) begin
        mem_7 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_8 <= 32'hb52023;
    end else begin
      if (11'h8 == _T_12323) begin
        mem_8 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_9 <= 32'hb52023;
    end else begin
      if (11'h9 == _T_12323) begin
        mem_9 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_10 <= 32'h7400593;
    end else begin
      if (11'ha == _T_12323) begin
        mem_10 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_11 <= 32'hb52023;
    end else begin
      if (11'hb == _T_12323) begin
        mem_11 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_12 <= 32'h6500593;
    end else begin
      if (11'hc == _T_12323) begin
        mem_12 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_13 <= 32'hb52023;
    end else begin
      if (11'hd == _T_12323) begin
        mem_13 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_14 <= 32'h6400593;
    end else begin
      if (11'he == _T_12323) begin
        mem_14 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_15 <= 32'hb52023;
    end else begin
      if (11'hf == _T_12323) begin
        mem_15 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_16 <= 32'h2100593;
    end else begin
      if (11'h10 == _T_12323) begin
        mem_16 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_17 <= 32'hb52023;
    end else begin
      if (11'h11 == _T_12323) begin
        mem_17 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_18 <= 32'ha00593;
    end else begin
      if (11'h12 == _T_12323) begin
        mem_18 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_19 <= 32'hb52023;
    end else begin
      if (11'h13 == _T_12323) begin
        mem_19 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_20 <= 32'h0;
    end else begin
      if (11'h14 == _T_12323) begin
        mem_20 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_21 <= 32'h0;
    end else begin
      if (11'h15 == _T_12323) begin
        mem_21 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_22 <= 32'h0;
    end else begin
      if (11'h16 == _T_12323) begin
        mem_22 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_23 <= 32'h0;
    end else begin
      if (11'h17 == _T_12323) begin
        mem_23 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_24 <= 32'h0;
    end else begin
      if (11'h18 == _T_12323) begin
        mem_24 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_25 <= 32'h0;
    end else begin
      if (11'h19 == _T_12323) begin
        mem_25 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_26 <= 32'h0;
    end else begin
      if (11'h1a == _T_12323) begin
        mem_26 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_27 <= 32'h0;
    end else begin
      if (11'h1b == _T_12323) begin
        mem_27 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_28 <= 32'h0;
    end else begin
      if (11'h1c == _T_12323) begin
        mem_28 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_29 <= 32'h0;
    end else begin
      if (11'h1d == _T_12323) begin
        mem_29 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_30 <= 32'h0;
    end else begin
      if (11'h1e == _T_12323) begin
        mem_30 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_31 <= 32'h0;
    end else begin
      if (11'h1f == _T_12323) begin
        mem_31 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_32 <= 32'h0;
    end else begin
      if (11'h20 == _T_12323) begin
        mem_32 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_33 <= 32'h0;
    end else begin
      if (11'h21 == _T_12323) begin
        mem_33 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_34 <= 32'h0;
    end else begin
      if (11'h22 == _T_12323) begin
        mem_34 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_35 <= 32'h0;
    end else begin
      if (11'h23 == _T_12323) begin
        mem_35 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_36 <= 32'h0;
    end else begin
      if (11'h24 == _T_12323) begin
        mem_36 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_37 <= 32'h0;
    end else begin
      if (11'h25 == _T_12323) begin
        mem_37 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_38 <= 32'h0;
    end else begin
      if (11'h26 == _T_12323) begin
        mem_38 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_39 <= 32'h0;
    end else begin
      if (11'h27 == _T_12323) begin
        mem_39 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_40 <= 32'h0;
    end else begin
      if (11'h28 == _T_12323) begin
        mem_40 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_41 <= 32'h0;
    end else begin
      if (11'h29 == _T_12323) begin
        mem_41 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_42 <= 32'h0;
    end else begin
      if (11'h2a == _T_12323) begin
        mem_42 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_43 <= 32'h0;
    end else begin
      if (11'h2b == _T_12323) begin
        mem_43 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_44 <= 32'h0;
    end else begin
      if (11'h2c == _T_12323) begin
        mem_44 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_45 <= 32'h0;
    end else begin
      if (11'h2d == _T_12323) begin
        mem_45 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_46 <= 32'h0;
    end else begin
      if (11'h2e == _T_12323) begin
        mem_46 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_47 <= 32'h0;
    end else begin
      if (11'h2f == _T_12323) begin
        mem_47 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_48 <= 32'h0;
    end else begin
      if (11'h30 == _T_12323) begin
        mem_48 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_49 <= 32'h0;
    end else begin
      if (11'h31 == _T_12323) begin
        mem_49 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_50 <= 32'h0;
    end else begin
      if (11'h32 == _T_12323) begin
        mem_50 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_51 <= 32'h0;
    end else begin
      if (11'h33 == _T_12323) begin
        mem_51 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_52 <= 32'h0;
    end else begin
      if (11'h34 == _T_12323) begin
        mem_52 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_53 <= 32'h0;
    end else begin
      if (11'h35 == _T_12323) begin
        mem_53 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_54 <= 32'h0;
    end else begin
      if (11'h36 == _T_12323) begin
        mem_54 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_55 <= 32'h0;
    end else begin
      if (11'h37 == _T_12323) begin
        mem_55 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_56 <= 32'h0;
    end else begin
      if (11'h38 == _T_12323) begin
        mem_56 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_57 <= 32'h0;
    end else begin
      if (11'h39 == _T_12323) begin
        mem_57 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_58 <= 32'h0;
    end else begin
      if (11'h3a == _T_12323) begin
        mem_58 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_59 <= 32'h0;
    end else begin
      if (11'h3b == _T_12323) begin
        mem_59 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_60 <= 32'h0;
    end else begin
      if (11'h3c == _T_12323) begin
        mem_60 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_61 <= 32'h0;
    end else begin
      if (11'h3d == _T_12323) begin
        mem_61 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_62 <= 32'h0;
    end else begin
      if (11'h3e == _T_12323) begin
        mem_62 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_63 <= 32'h0;
    end else begin
      if (11'h3f == _T_12323) begin
        mem_63 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_64 <= 32'h0;
    end else begin
      if (11'h40 == _T_12323) begin
        mem_64 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_65 <= 32'h0;
    end else begin
      if (11'h41 == _T_12323) begin
        mem_65 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_66 <= 32'h0;
    end else begin
      if (11'h42 == _T_12323) begin
        mem_66 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_67 <= 32'h0;
    end else begin
      if (11'h43 == _T_12323) begin
        mem_67 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_68 <= 32'h0;
    end else begin
      if (11'h44 == _T_12323) begin
        mem_68 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_69 <= 32'h0;
    end else begin
      if (11'h45 == _T_12323) begin
        mem_69 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_70 <= 32'h0;
    end else begin
      if (11'h46 == _T_12323) begin
        mem_70 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_71 <= 32'h0;
    end else begin
      if (11'h47 == _T_12323) begin
        mem_71 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_72 <= 32'h0;
    end else begin
      if (11'h48 == _T_12323) begin
        mem_72 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_73 <= 32'h0;
    end else begin
      if (11'h49 == _T_12323) begin
        mem_73 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_74 <= 32'h0;
    end else begin
      if (11'h4a == _T_12323) begin
        mem_74 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_75 <= 32'h0;
    end else begin
      if (11'h4b == _T_12323) begin
        mem_75 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_76 <= 32'h0;
    end else begin
      if (11'h4c == _T_12323) begin
        mem_76 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_77 <= 32'h0;
    end else begin
      if (11'h4d == _T_12323) begin
        mem_77 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_78 <= 32'h0;
    end else begin
      if (11'h4e == _T_12323) begin
        mem_78 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_79 <= 32'h0;
    end else begin
      if (11'h4f == _T_12323) begin
        mem_79 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_80 <= 32'h0;
    end else begin
      if (11'h50 == _T_12323) begin
        mem_80 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_81 <= 32'h0;
    end else begin
      if (11'h51 == _T_12323) begin
        mem_81 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_82 <= 32'h0;
    end else begin
      if (11'h52 == _T_12323) begin
        mem_82 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_83 <= 32'h0;
    end else begin
      if (11'h53 == _T_12323) begin
        mem_83 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_84 <= 32'h0;
    end else begin
      if (11'h54 == _T_12323) begin
        mem_84 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_85 <= 32'h0;
    end else begin
      if (11'h55 == _T_12323) begin
        mem_85 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_86 <= 32'h0;
    end else begin
      if (11'h56 == _T_12323) begin
        mem_86 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_87 <= 32'h0;
    end else begin
      if (11'h57 == _T_12323) begin
        mem_87 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_88 <= 32'h0;
    end else begin
      if (11'h58 == _T_12323) begin
        mem_88 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_89 <= 32'h0;
    end else begin
      if (11'h59 == _T_12323) begin
        mem_89 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_90 <= 32'h0;
    end else begin
      if (11'h5a == _T_12323) begin
        mem_90 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_91 <= 32'h0;
    end else begin
      if (11'h5b == _T_12323) begin
        mem_91 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_92 <= 32'h0;
    end else begin
      if (11'h5c == _T_12323) begin
        mem_92 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_93 <= 32'h0;
    end else begin
      if (11'h5d == _T_12323) begin
        mem_93 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_94 <= 32'h0;
    end else begin
      if (11'h5e == _T_12323) begin
        mem_94 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_95 <= 32'h0;
    end else begin
      if (11'h5f == _T_12323) begin
        mem_95 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_96 <= 32'h0;
    end else begin
      if (11'h60 == _T_12323) begin
        mem_96 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_97 <= 32'h0;
    end else begin
      if (11'h61 == _T_12323) begin
        mem_97 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_98 <= 32'h0;
    end else begin
      if (11'h62 == _T_12323) begin
        mem_98 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_99 <= 32'h0;
    end else begin
      if (11'h63 == _T_12323) begin
        mem_99 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_100 <= 32'h0;
    end else begin
      if (11'h64 == _T_12323) begin
        mem_100 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_101 <= 32'h0;
    end else begin
      if (11'h65 == _T_12323) begin
        mem_101 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_102 <= 32'h0;
    end else begin
      if (11'h66 == _T_12323) begin
        mem_102 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_103 <= 32'h0;
    end else begin
      if (11'h67 == _T_12323) begin
        mem_103 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_104 <= 32'h0;
    end else begin
      if (11'h68 == _T_12323) begin
        mem_104 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_105 <= 32'h0;
    end else begin
      if (11'h69 == _T_12323) begin
        mem_105 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_106 <= 32'h0;
    end else begin
      if (11'h6a == _T_12323) begin
        mem_106 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_107 <= 32'h0;
    end else begin
      if (11'h6b == _T_12323) begin
        mem_107 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_108 <= 32'h0;
    end else begin
      if (11'h6c == _T_12323) begin
        mem_108 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_109 <= 32'h0;
    end else begin
      if (11'h6d == _T_12323) begin
        mem_109 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_110 <= 32'h0;
    end else begin
      if (11'h6e == _T_12323) begin
        mem_110 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_111 <= 32'h0;
    end else begin
      if (11'h6f == _T_12323) begin
        mem_111 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_112 <= 32'h0;
    end else begin
      if (11'h70 == _T_12323) begin
        mem_112 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_113 <= 32'h0;
    end else begin
      if (11'h71 == _T_12323) begin
        mem_113 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_114 <= 32'h0;
    end else begin
      if (11'h72 == _T_12323) begin
        mem_114 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_115 <= 32'h0;
    end else begin
      if (11'h73 == _T_12323) begin
        mem_115 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_116 <= 32'h0;
    end else begin
      if (11'h74 == _T_12323) begin
        mem_116 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_117 <= 32'h0;
    end else begin
      if (11'h75 == _T_12323) begin
        mem_117 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_118 <= 32'h0;
    end else begin
      if (11'h76 == _T_12323) begin
        mem_118 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_119 <= 32'h0;
    end else begin
      if (11'h77 == _T_12323) begin
        mem_119 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_120 <= 32'h0;
    end else begin
      if (11'h78 == _T_12323) begin
        mem_120 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_121 <= 32'h0;
    end else begin
      if (11'h79 == _T_12323) begin
        mem_121 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_122 <= 32'h0;
    end else begin
      if (11'h7a == _T_12323) begin
        mem_122 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_123 <= 32'h0;
    end else begin
      if (11'h7b == _T_12323) begin
        mem_123 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_124 <= 32'h0;
    end else begin
      if (11'h7c == _T_12323) begin
        mem_124 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_125 <= 32'h0;
    end else begin
      if (11'h7d == _T_12323) begin
        mem_125 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_126 <= 32'h0;
    end else begin
      if (11'h7e == _T_12323) begin
        mem_126 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_127 <= 32'h0;
    end else begin
      if (11'h7f == _T_12323) begin
        mem_127 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_128 <= 32'h0;
    end else begin
      if (11'h80 == _T_12323) begin
        mem_128 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_129 <= 32'h0;
    end else begin
      if (11'h81 == _T_12323) begin
        mem_129 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_130 <= 32'h0;
    end else begin
      if (11'h82 == _T_12323) begin
        mem_130 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_131 <= 32'h0;
    end else begin
      if (11'h83 == _T_12323) begin
        mem_131 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_132 <= 32'h0;
    end else begin
      if (11'h84 == _T_12323) begin
        mem_132 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_133 <= 32'h0;
    end else begin
      if (11'h85 == _T_12323) begin
        mem_133 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_134 <= 32'h0;
    end else begin
      if (11'h86 == _T_12323) begin
        mem_134 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_135 <= 32'h0;
    end else begin
      if (11'h87 == _T_12323) begin
        mem_135 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_136 <= 32'h0;
    end else begin
      if (11'h88 == _T_12323) begin
        mem_136 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_137 <= 32'h0;
    end else begin
      if (11'h89 == _T_12323) begin
        mem_137 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_138 <= 32'h0;
    end else begin
      if (11'h8a == _T_12323) begin
        mem_138 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_139 <= 32'h0;
    end else begin
      if (11'h8b == _T_12323) begin
        mem_139 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_140 <= 32'h0;
    end else begin
      if (11'h8c == _T_12323) begin
        mem_140 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_141 <= 32'h0;
    end else begin
      if (11'h8d == _T_12323) begin
        mem_141 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_142 <= 32'h0;
    end else begin
      if (11'h8e == _T_12323) begin
        mem_142 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_143 <= 32'h0;
    end else begin
      if (11'h8f == _T_12323) begin
        mem_143 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_144 <= 32'h0;
    end else begin
      if (11'h90 == _T_12323) begin
        mem_144 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_145 <= 32'h0;
    end else begin
      if (11'h91 == _T_12323) begin
        mem_145 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_146 <= 32'h0;
    end else begin
      if (11'h92 == _T_12323) begin
        mem_146 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_147 <= 32'h0;
    end else begin
      if (11'h93 == _T_12323) begin
        mem_147 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_148 <= 32'h0;
    end else begin
      if (11'h94 == _T_12323) begin
        mem_148 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_149 <= 32'h0;
    end else begin
      if (11'h95 == _T_12323) begin
        mem_149 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_150 <= 32'h0;
    end else begin
      if (11'h96 == _T_12323) begin
        mem_150 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_151 <= 32'h0;
    end else begin
      if (11'h97 == _T_12323) begin
        mem_151 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_152 <= 32'h0;
    end else begin
      if (11'h98 == _T_12323) begin
        mem_152 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_153 <= 32'h0;
    end else begin
      if (11'h99 == _T_12323) begin
        mem_153 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_154 <= 32'h0;
    end else begin
      if (11'h9a == _T_12323) begin
        mem_154 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_155 <= 32'h0;
    end else begin
      if (11'h9b == _T_12323) begin
        mem_155 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_156 <= 32'h0;
    end else begin
      if (11'h9c == _T_12323) begin
        mem_156 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_157 <= 32'h0;
    end else begin
      if (11'h9d == _T_12323) begin
        mem_157 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_158 <= 32'h0;
    end else begin
      if (11'h9e == _T_12323) begin
        mem_158 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_159 <= 32'h0;
    end else begin
      if (11'h9f == _T_12323) begin
        mem_159 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_160 <= 32'h0;
    end else begin
      if (11'ha0 == _T_12323) begin
        mem_160 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_161 <= 32'h0;
    end else begin
      if (11'ha1 == _T_12323) begin
        mem_161 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_162 <= 32'h0;
    end else begin
      if (11'ha2 == _T_12323) begin
        mem_162 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_163 <= 32'h0;
    end else begin
      if (11'ha3 == _T_12323) begin
        mem_163 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_164 <= 32'h0;
    end else begin
      if (11'ha4 == _T_12323) begin
        mem_164 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_165 <= 32'h0;
    end else begin
      if (11'ha5 == _T_12323) begin
        mem_165 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_166 <= 32'h0;
    end else begin
      if (11'ha6 == _T_12323) begin
        mem_166 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_167 <= 32'h0;
    end else begin
      if (11'ha7 == _T_12323) begin
        mem_167 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_168 <= 32'h0;
    end else begin
      if (11'ha8 == _T_12323) begin
        mem_168 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_169 <= 32'h0;
    end else begin
      if (11'ha9 == _T_12323) begin
        mem_169 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_170 <= 32'h0;
    end else begin
      if (11'haa == _T_12323) begin
        mem_170 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_171 <= 32'h0;
    end else begin
      if (11'hab == _T_12323) begin
        mem_171 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_172 <= 32'h0;
    end else begin
      if (11'hac == _T_12323) begin
        mem_172 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_173 <= 32'h0;
    end else begin
      if (11'had == _T_12323) begin
        mem_173 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_174 <= 32'h0;
    end else begin
      if (11'hae == _T_12323) begin
        mem_174 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_175 <= 32'h0;
    end else begin
      if (11'haf == _T_12323) begin
        mem_175 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_176 <= 32'h0;
    end else begin
      if (11'hb0 == _T_12323) begin
        mem_176 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_177 <= 32'h0;
    end else begin
      if (11'hb1 == _T_12323) begin
        mem_177 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_178 <= 32'h0;
    end else begin
      if (11'hb2 == _T_12323) begin
        mem_178 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_179 <= 32'h0;
    end else begin
      if (11'hb3 == _T_12323) begin
        mem_179 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_180 <= 32'h0;
    end else begin
      if (11'hb4 == _T_12323) begin
        mem_180 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_181 <= 32'h0;
    end else begin
      if (11'hb5 == _T_12323) begin
        mem_181 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_182 <= 32'h0;
    end else begin
      if (11'hb6 == _T_12323) begin
        mem_182 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_183 <= 32'h0;
    end else begin
      if (11'hb7 == _T_12323) begin
        mem_183 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_184 <= 32'h0;
    end else begin
      if (11'hb8 == _T_12323) begin
        mem_184 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_185 <= 32'h0;
    end else begin
      if (11'hb9 == _T_12323) begin
        mem_185 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_186 <= 32'h0;
    end else begin
      if (11'hba == _T_12323) begin
        mem_186 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_187 <= 32'h0;
    end else begin
      if (11'hbb == _T_12323) begin
        mem_187 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_188 <= 32'h0;
    end else begin
      if (11'hbc == _T_12323) begin
        mem_188 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_189 <= 32'h0;
    end else begin
      if (11'hbd == _T_12323) begin
        mem_189 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_190 <= 32'h0;
    end else begin
      if (11'hbe == _T_12323) begin
        mem_190 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_191 <= 32'h0;
    end else begin
      if (11'hbf == _T_12323) begin
        mem_191 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_192 <= 32'h0;
    end else begin
      if (11'hc0 == _T_12323) begin
        mem_192 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_193 <= 32'h0;
    end else begin
      if (11'hc1 == _T_12323) begin
        mem_193 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_194 <= 32'h0;
    end else begin
      if (11'hc2 == _T_12323) begin
        mem_194 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_195 <= 32'h0;
    end else begin
      if (11'hc3 == _T_12323) begin
        mem_195 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_196 <= 32'h0;
    end else begin
      if (11'hc4 == _T_12323) begin
        mem_196 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_197 <= 32'h0;
    end else begin
      if (11'hc5 == _T_12323) begin
        mem_197 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_198 <= 32'h0;
    end else begin
      if (11'hc6 == _T_12323) begin
        mem_198 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_199 <= 32'h0;
    end else begin
      if (11'hc7 == _T_12323) begin
        mem_199 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_200 <= 32'h0;
    end else begin
      if (11'hc8 == _T_12323) begin
        mem_200 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_201 <= 32'h0;
    end else begin
      if (11'hc9 == _T_12323) begin
        mem_201 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_202 <= 32'h0;
    end else begin
      if (11'hca == _T_12323) begin
        mem_202 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_203 <= 32'h0;
    end else begin
      if (11'hcb == _T_12323) begin
        mem_203 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_204 <= 32'h0;
    end else begin
      if (11'hcc == _T_12323) begin
        mem_204 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_205 <= 32'h0;
    end else begin
      if (11'hcd == _T_12323) begin
        mem_205 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_206 <= 32'h0;
    end else begin
      if (11'hce == _T_12323) begin
        mem_206 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_207 <= 32'h0;
    end else begin
      if (11'hcf == _T_12323) begin
        mem_207 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_208 <= 32'h0;
    end else begin
      if (11'hd0 == _T_12323) begin
        mem_208 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_209 <= 32'h0;
    end else begin
      if (11'hd1 == _T_12323) begin
        mem_209 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_210 <= 32'h0;
    end else begin
      if (11'hd2 == _T_12323) begin
        mem_210 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_211 <= 32'h0;
    end else begin
      if (11'hd3 == _T_12323) begin
        mem_211 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_212 <= 32'h0;
    end else begin
      if (11'hd4 == _T_12323) begin
        mem_212 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_213 <= 32'h0;
    end else begin
      if (11'hd5 == _T_12323) begin
        mem_213 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_214 <= 32'h0;
    end else begin
      if (11'hd6 == _T_12323) begin
        mem_214 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_215 <= 32'h0;
    end else begin
      if (11'hd7 == _T_12323) begin
        mem_215 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_216 <= 32'h0;
    end else begin
      if (11'hd8 == _T_12323) begin
        mem_216 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_217 <= 32'h0;
    end else begin
      if (11'hd9 == _T_12323) begin
        mem_217 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_218 <= 32'h0;
    end else begin
      if (11'hda == _T_12323) begin
        mem_218 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_219 <= 32'h0;
    end else begin
      if (11'hdb == _T_12323) begin
        mem_219 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_220 <= 32'h0;
    end else begin
      if (11'hdc == _T_12323) begin
        mem_220 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_221 <= 32'h0;
    end else begin
      if (11'hdd == _T_12323) begin
        mem_221 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_222 <= 32'h0;
    end else begin
      if (11'hde == _T_12323) begin
        mem_222 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_223 <= 32'h0;
    end else begin
      if (11'hdf == _T_12323) begin
        mem_223 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_224 <= 32'h0;
    end else begin
      if (11'he0 == _T_12323) begin
        mem_224 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_225 <= 32'h0;
    end else begin
      if (11'he1 == _T_12323) begin
        mem_225 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_226 <= 32'h0;
    end else begin
      if (11'he2 == _T_12323) begin
        mem_226 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_227 <= 32'h0;
    end else begin
      if (11'he3 == _T_12323) begin
        mem_227 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_228 <= 32'h0;
    end else begin
      if (11'he4 == _T_12323) begin
        mem_228 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_229 <= 32'h0;
    end else begin
      if (11'he5 == _T_12323) begin
        mem_229 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_230 <= 32'h0;
    end else begin
      if (11'he6 == _T_12323) begin
        mem_230 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_231 <= 32'h0;
    end else begin
      if (11'he7 == _T_12323) begin
        mem_231 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_232 <= 32'h0;
    end else begin
      if (11'he8 == _T_12323) begin
        mem_232 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_233 <= 32'h0;
    end else begin
      if (11'he9 == _T_12323) begin
        mem_233 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_234 <= 32'h0;
    end else begin
      if (11'hea == _T_12323) begin
        mem_234 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_235 <= 32'h0;
    end else begin
      if (11'heb == _T_12323) begin
        mem_235 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_236 <= 32'h0;
    end else begin
      if (11'hec == _T_12323) begin
        mem_236 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_237 <= 32'h0;
    end else begin
      if (11'hed == _T_12323) begin
        mem_237 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_238 <= 32'h0;
    end else begin
      if (11'hee == _T_12323) begin
        mem_238 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_239 <= 32'h0;
    end else begin
      if (11'hef == _T_12323) begin
        mem_239 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_240 <= 32'h0;
    end else begin
      if (11'hf0 == _T_12323) begin
        mem_240 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_241 <= 32'h0;
    end else begin
      if (11'hf1 == _T_12323) begin
        mem_241 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_242 <= 32'h0;
    end else begin
      if (11'hf2 == _T_12323) begin
        mem_242 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_243 <= 32'h0;
    end else begin
      if (11'hf3 == _T_12323) begin
        mem_243 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_244 <= 32'h0;
    end else begin
      if (11'hf4 == _T_12323) begin
        mem_244 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_245 <= 32'h0;
    end else begin
      if (11'hf5 == _T_12323) begin
        mem_245 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_246 <= 32'h0;
    end else begin
      if (11'hf6 == _T_12323) begin
        mem_246 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_247 <= 32'h0;
    end else begin
      if (11'hf7 == _T_12323) begin
        mem_247 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_248 <= 32'h0;
    end else begin
      if (11'hf8 == _T_12323) begin
        mem_248 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_249 <= 32'h0;
    end else begin
      if (11'hf9 == _T_12323) begin
        mem_249 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_250 <= 32'h0;
    end else begin
      if (11'hfa == _T_12323) begin
        mem_250 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_251 <= 32'h0;
    end else begin
      if (11'hfb == _T_12323) begin
        mem_251 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_252 <= 32'h0;
    end else begin
      if (11'hfc == _T_12323) begin
        mem_252 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_253 <= 32'h0;
    end else begin
      if (11'hfd == _T_12323) begin
        mem_253 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_254 <= 32'h0;
    end else begin
      if (11'hfe == _T_12323) begin
        mem_254 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_255 <= 32'h0;
    end else begin
      if (11'hff == _T_12323) begin
        mem_255 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_256 <= 32'h0;
    end else begin
      if (11'h100 == _T_12323) begin
        mem_256 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_257 <= 32'h0;
    end else begin
      if (11'h101 == _T_12323) begin
        mem_257 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_258 <= 32'h0;
    end else begin
      if (11'h102 == _T_12323) begin
        mem_258 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_259 <= 32'h0;
    end else begin
      if (11'h103 == _T_12323) begin
        mem_259 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_260 <= 32'h0;
    end else begin
      if (11'h104 == _T_12323) begin
        mem_260 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_261 <= 32'h0;
    end else begin
      if (11'h105 == _T_12323) begin
        mem_261 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_262 <= 32'h0;
    end else begin
      if (11'h106 == _T_12323) begin
        mem_262 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_263 <= 32'h0;
    end else begin
      if (11'h107 == _T_12323) begin
        mem_263 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_264 <= 32'h0;
    end else begin
      if (11'h108 == _T_12323) begin
        mem_264 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_265 <= 32'h0;
    end else begin
      if (11'h109 == _T_12323) begin
        mem_265 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_266 <= 32'h0;
    end else begin
      if (11'h10a == _T_12323) begin
        mem_266 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_267 <= 32'h0;
    end else begin
      if (11'h10b == _T_12323) begin
        mem_267 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_268 <= 32'h0;
    end else begin
      if (11'h10c == _T_12323) begin
        mem_268 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_269 <= 32'h0;
    end else begin
      if (11'h10d == _T_12323) begin
        mem_269 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_270 <= 32'h0;
    end else begin
      if (11'h10e == _T_12323) begin
        mem_270 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_271 <= 32'h0;
    end else begin
      if (11'h10f == _T_12323) begin
        mem_271 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_272 <= 32'h0;
    end else begin
      if (11'h110 == _T_12323) begin
        mem_272 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_273 <= 32'h0;
    end else begin
      if (11'h111 == _T_12323) begin
        mem_273 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_274 <= 32'h0;
    end else begin
      if (11'h112 == _T_12323) begin
        mem_274 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_275 <= 32'h0;
    end else begin
      if (11'h113 == _T_12323) begin
        mem_275 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_276 <= 32'h0;
    end else begin
      if (11'h114 == _T_12323) begin
        mem_276 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_277 <= 32'h0;
    end else begin
      if (11'h115 == _T_12323) begin
        mem_277 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_278 <= 32'h0;
    end else begin
      if (11'h116 == _T_12323) begin
        mem_278 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_279 <= 32'h0;
    end else begin
      if (11'h117 == _T_12323) begin
        mem_279 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_280 <= 32'h0;
    end else begin
      if (11'h118 == _T_12323) begin
        mem_280 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_281 <= 32'h0;
    end else begin
      if (11'h119 == _T_12323) begin
        mem_281 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_282 <= 32'h0;
    end else begin
      if (11'h11a == _T_12323) begin
        mem_282 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_283 <= 32'h0;
    end else begin
      if (11'h11b == _T_12323) begin
        mem_283 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_284 <= 32'h0;
    end else begin
      if (11'h11c == _T_12323) begin
        mem_284 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_285 <= 32'h0;
    end else begin
      if (11'h11d == _T_12323) begin
        mem_285 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_286 <= 32'h0;
    end else begin
      if (11'h11e == _T_12323) begin
        mem_286 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_287 <= 32'h0;
    end else begin
      if (11'h11f == _T_12323) begin
        mem_287 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_288 <= 32'h0;
    end else begin
      if (11'h120 == _T_12323) begin
        mem_288 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_289 <= 32'h0;
    end else begin
      if (11'h121 == _T_12323) begin
        mem_289 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_290 <= 32'h0;
    end else begin
      if (11'h122 == _T_12323) begin
        mem_290 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_291 <= 32'h0;
    end else begin
      if (11'h123 == _T_12323) begin
        mem_291 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_292 <= 32'h0;
    end else begin
      if (11'h124 == _T_12323) begin
        mem_292 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_293 <= 32'h0;
    end else begin
      if (11'h125 == _T_12323) begin
        mem_293 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_294 <= 32'h0;
    end else begin
      if (11'h126 == _T_12323) begin
        mem_294 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_295 <= 32'h0;
    end else begin
      if (11'h127 == _T_12323) begin
        mem_295 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_296 <= 32'h0;
    end else begin
      if (11'h128 == _T_12323) begin
        mem_296 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_297 <= 32'h0;
    end else begin
      if (11'h129 == _T_12323) begin
        mem_297 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_298 <= 32'h0;
    end else begin
      if (11'h12a == _T_12323) begin
        mem_298 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_299 <= 32'h0;
    end else begin
      if (11'h12b == _T_12323) begin
        mem_299 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_300 <= 32'h0;
    end else begin
      if (11'h12c == _T_12323) begin
        mem_300 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_301 <= 32'h0;
    end else begin
      if (11'h12d == _T_12323) begin
        mem_301 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_302 <= 32'h0;
    end else begin
      if (11'h12e == _T_12323) begin
        mem_302 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_303 <= 32'h0;
    end else begin
      if (11'h12f == _T_12323) begin
        mem_303 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_304 <= 32'h0;
    end else begin
      if (11'h130 == _T_12323) begin
        mem_304 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_305 <= 32'h0;
    end else begin
      if (11'h131 == _T_12323) begin
        mem_305 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_306 <= 32'h0;
    end else begin
      if (11'h132 == _T_12323) begin
        mem_306 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_307 <= 32'h0;
    end else begin
      if (11'h133 == _T_12323) begin
        mem_307 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_308 <= 32'h0;
    end else begin
      if (11'h134 == _T_12323) begin
        mem_308 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_309 <= 32'h0;
    end else begin
      if (11'h135 == _T_12323) begin
        mem_309 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_310 <= 32'h0;
    end else begin
      if (11'h136 == _T_12323) begin
        mem_310 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_311 <= 32'h0;
    end else begin
      if (11'h137 == _T_12323) begin
        mem_311 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_312 <= 32'h0;
    end else begin
      if (11'h138 == _T_12323) begin
        mem_312 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_313 <= 32'h0;
    end else begin
      if (11'h139 == _T_12323) begin
        mem_313 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_314 <= 32'h0;
    end else begin
      if (11'h13a == _T_12323) begin
        mem_314 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_315 <= 32'h0;
    end else begin
      if (11'h13b == _T_12323) begin
        mem_315 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_316 <= 32'h0;
    end else begin
      if (11'h13c == _T_12323) begin
        mem_316 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_317 <= 32'h0;
    end else begin
      if (11'h13d == _T_12323) begin
        mem_317 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_318 <= 32'h0;
    end else begin
      if (11'h13e == _T_12323) begin
        mem_318 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_319 <= 32'h0;
    end else begin
      if (11'h13f == _T_12323) begin
        mem_319 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_320 <= 32'h0;
    end else begin
      if (11'h140 == _T_12323) begin
        mem_320 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_321 <= 32'h0;
    end else begin
      if (11'h141 == _T_12323) begin
        mem_321 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_322 <= 32'h0;
    end else begin
      if (11'h142 == _T_12323) begin
        mem_322 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_323 <= 32'h0;
    end else begin
      if (11'h143 == _T_12323) begin
        mem_323 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_324 <= 32'h0;
    end else begin
      if (11'h144 == _T_12323) begin
        mem_324 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_325 <= 32'h0;
    end else begin
      if (11'h145 == _T_12323) begin
        mem_325 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_326 <= 32'h0;
    end else begin
      if (11'h146 == _T_12323) begin
        mem_326 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_327 <= 32'h0;
    end else begin
      if (11'h147 == _T_12323) begin
        mem_327 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_328 <= 32'h0;
    end else begin
      if (11'h148 == _T_12323) begin
        mem_328 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_329 <= 32'h0;
    end else begin
      if (11'h149 == _T_12323) begin
        mem_329 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_330 <= 32'h0;
    end else begin
      if (11'h14a == _T_12323) begin
        mem_330 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_331 <= 32'h0;
    end else begin
      if (11'h14b == _T_12323) begin
        mem_331 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_332 <= 32'h0;
    end else begin
      if (11'h14c == _T_12323) begin
        mem_332 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_333 <= 32'h0;
    end else begin
      if (11'h14d == _T_12323) begin
        mem_333 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_334 <= 32'h0;
    end else begin
      if (11'h14e == _T_12323) begin
        mem_334 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_335 <= 32'h0;
    end else begin
      if (11'h14f == _T_12323) begin
        mem_335 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_336 <= 32'h0;
    end else begin
      if (11'h150 == _T_12323) begin
        mem_336 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_337 <= 32'h0;
    end else begin
      if (11'h151 == _T_12323) begin
        mem_337 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_338 <= 32'h0;
    end else begin
      if (11'h152 == _T_12323) begin
        mem_338 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_339 <= 32'h0;
    end else begin
      if (11'h153 == _T_12323) begin
        mem_339 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_340 <= 32'h0;
    end else begin
      if (11'h154 == _T_12323) begin
        mem_340 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_341 <= 32'h0;
    end else begin
      if (11'h155 == _T_12323) begin
        mem_341 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_342 <= 32'h0;
    end else begin
      if (11'h156 == _T_12323) begin
        mem_342 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_343 <= 32'h0;
    end else begin
      if (11'h157 == _T_12323) begin
        mem_343 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_344 <= 32'h0;
    end else begin
      if (11'h158 == _T_12323) begin
        mem_344 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_345 <= 32'h0;
    end else begin
      if (11'h159 == _T_12323) begin
        mem_345 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_346 <= 32'h0;
    end else begin
      if (11'h15a == _T_12323) begin
        mem_346 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_347 <= 32'h0;
    end else begin
      if (11'h15b == _T_12323) begin
        mem_347 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_348 <= 32'h0;
    end else begin
      if (11'h15c == _T_12323) begin
        mem_348 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_349 <= 32'h0;
    end else begin
      if (11'h15d == _T_12323) begin
        mem_349 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_350 <= 32'h0;
    end else begin
      if (11'h15e == _T_12323) begin
        mem_350 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_351 <= 32'h0;
    end else begin
      if (11'h15f == _T_12323) begin
        mem_351 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_352 <= 32'h0;
    end else begin
      if (11'h160 == _T_12323) begin
        mem_352 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_353 <= 32'h0;
    end else begin
      if (11'h161 == _T_12323) begin
        mem_353 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_354 <= 32'h0;
    end else begin
      if (11'h162 == _T_12323) begin
        mem_354 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_355 <= 32'h0;
    end else begin
      if (11'h163 == _T_12323) begin
        mem_355 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_356 <= 32'h0;
    end else begin
      if (11'h164 == _T_12323) begin
        mem_356 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_357 <= 32'h0;
    end else begin
      if (11'h165 == _T_12323) begin
        mem_357 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_358 <= 32'h0;
    end else begin
      if (11'h166 == _T_12323) begin
        mem_358 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_359 <= 32'h0;
    end else begin
      if (11'h167 == _T_12323) begin
        mem_359 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_360 <= 32'h0;
    end else begin
      if (11'h168 == _T_12323) begin
        mem_360 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_361 <= 32'h0;
    end else begin
      if (11'h169 == _T_12323) begin
        mem_361 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_362 <= 32'h0;
    end else begin
      if (11'h16a == _T_12323) begin
        mem_362 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_363 <= 32'h0;
    end else begin
      if (11'h16b == _T_12323) begin
        mem_363 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_364 <= 32'h0;
    end else begin
      if (11'h16c == _T_12323) begin
        mem_364 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_365 <= 32'h0;
    end else begin
      if (11'h16d == _T_12323) begin
        mem_365 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_366 <= 32'h0;
    end else begin
      if (11'h16e == _T_12323) begin
        mem_366 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_367 <= 32'h0;
    end else begin
      if (11'h16f == _T_12323) begin
        mem_367 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_368 <= 32'h0;
    end else begin
      if (11'h170 == _T_12323) begin
        mem_368 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_369 <= 32'h0;
    end else begin
      if (11'h171 == _T_12323) begin
        mem_369 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_370 <= 32'h0;
    end else begin
      if (11'h172 == _T_12323) begin
        mem_370 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_371 <= 32'h0;
    end else begin
      if (11'h173 == _T_12323) begin
        mem_371 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_372 <= 32'h0;
    end else begin
      if (11'h174 == _T_12323) begin
        mem_372 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_373 <= 32'h0;
    end else begin
      if (11'h175 == _T_12323) begin
        mem_373 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_374 <= 32'h0;
    end else begin
      if (11'h176 == _T_12323) begin
        mem_374 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_375 <= 32'h0;
    end else begin
      if (11'h177 == _T_12323) begin
        mem_375 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_376 <= 32'h0;
    end else begin
      if (11'h178 == _T_12323) begin
        mem_376 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_377 <= 32'h0;
    end else begin
      if (11'h179 == _T_12323) begin
        mem_377 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_378 <= 32'h0;
    end else begin
      if (11'h17a == _T_12323) begin
        mem_378 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_379 <= 32'h0;
    end else begin
      if (11'h17b == _T_12323) begin
        mem_379 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_380 <= 32'h0;
    end else begin
      if (11'h17c == _T_12323) begin
        mem_380 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_381 <= 32'h0;
    end else begin
      if (11'h17d == _T_12323) begin
        mem_381 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_382 <= 32'h0;
    end else begin
      if (11'h17e == _T_12323) begin
        mem_382 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_383 <= 32'h0;
    end else begin
      if (11'h17f == _T_12323) begin
        mem_383 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_384 <= 32'h0;
    end else begin
      if (11'h180 == _T_12323) begin
        mem_384 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_385 <= 32'h0;
    end else begin
      if (11'h181 == _T_12323) begin
        mem_385 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_386 <= 32'h0;
    end else begin
      if (11'h182 == _T_12323) begin
        mem_386 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_387 <= 32'h0;
    end else begin
      if (11'h183 == _T_12323) begin
        mem_387 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_388 <= 32'h0;
    end else begin
      if (11'h184 == _T_12323) begin
        mem_388 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_389 <= 32'h0;
    end else begin
      if (11'h185 == _T_12323) begin
        mem_389 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_390 <= 32'h0;
    end else begin
      if (11'h186 == _T_12323) begin
        mem_390 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_391 <= 32'h0;
    end else begin
      if (11'h187 == _T_12323) begin
        mem_391 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_392 <= 32'h0;
    end else begin
      if (11'h188 == _T_12323) begin
        mem_392 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_393 <= 32'h0;
    end else begin
      if (11'h189 == _T_12323) begin
        mem_393 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_394 <= 32'h0;
    end else begin
      if (11'h18a == _T_12323) begin
        mem_394 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_395 <= 32'h0;
    end else begin
      if (11'h18b == _T_12323) begin
        mem_395 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_396 <= 32'h0;
    end else begin
      if (11'h18c == _T_12323) begin
        mem_396 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_397 <= 32'h0;
    end else begin
      if (11'h18d == _T_12323) begin
        mem_397 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_398 <= 32'h0;
    end else begin
      if (11'h18e == _T_12323) begin
        mem_398 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_399 <= 32'h0;
    end else begin
      if (11'h18f == _T_12323) begin
        mem_399 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_400 <= 32'h0;
    end else begin
      if (11'h190 == _T_12323) begin
        mem_400 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_401 <= 32'h0;
    end else begin
      if (11'h191 == _T_12323) begin
        mem_401 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_402 <= 32'h0;
    end else begin
      if (11'h192 == _T_12323) begin
        mem_402 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_403 <= 32'h0;
    end else begin
      if (11'h193 == _T_12323) begin
        mem_403 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_404 <= 32'h0;
    end else begin
      if (11'h194 == _T_12323) begin
        mem_404 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_405 <= 32'h0;
    end else begin
      if (11'h195 == _T_12323) begin
        mem_405 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_406 <= 32'h0;
    end else begin
      if (11'h196 == _T_12323) begin
        mem_406 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_407 <= 32'h0;
    end else begin
      if (11'h197 == _T_12323) begin
        mem_407 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_408 <= 32'h0;
    end else begin
      if (11'h198 == _T_12323) begin
        mem_408 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_409 <= 32'h0;
    end else begin
      if (11'h199 == _T_12323) begin
        mem_409 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_410 <= 32'h0;
    end else begin
      if (11'h19a == _T_12323) begin
        mem_410 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_411 <= 32'h0;
    end else begin
      if (11'h19b == _T_12323) begin
        mem_411 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_412 <= 32'h0;
    end else begin
      if (11'h19c == _T_12323) begin
        mem_412 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_413 <= 32'h0;
    end else begin
      if (11'h19d == _T_12323) begin
        mem_413 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_414 <= 32'h0;
    end else begin
      if (11'h19e == _T_12323) begin
        mem_414 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_415 <= 32'h0;
    end else begin
      if (11'h19f == _T_12323) begin
        mem_415 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_416 <= 32'h0;
    end else begin
      if (11'h1a0 == _T_12323) begin
        mem_416 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_417 <= 32'h0;
    end else begin
      if (11'h1a1 == _T_12323) begin
        mem_417 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_418 <= 32'h0;
    end else begin
      if (11'h1a2 == _T_12323) begin
        mem_418 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_419 <= 32'h0;
    end else begin
      if (11'h1a3 == _T_12323) begin
        mem_419 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_420 <= 32'h0;
    end else begin
      if (11'h1a4 == _T_12323) begin
        mem_420 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_421 <= 32'h0;
    end else begin
      if (11'h1a5 == _T_12323) begin
        mem_421 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_422 <= 32'h0;
    end else begin
      if (11'h1a6 == _T_12323) begin
        mem_422 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_423 <= 32'h0;
    end else begin
      if (11'h1a7 == _T_12323) begin
        mem_423 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_424 <= 32'h0;
    end else begin
      if (11'h1a8 == _T_12323) begin
        mem_424 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_425 <= 32'h0;
    end else begin
      if (11'h1a9 == _T_12323) begin
        mem_425 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_426 <= 32'h0;
    end else begin
      if (11'h1aa == _T_12323) begin
        mem_426 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_427 <= 32'h0;
    end else begin
      if (11'h1ab == _T_12323) begin
        mem_427 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_428 <= 32'h0;
    end else begin
      if (11'h1ac == _T_12323) begin
        mem_428 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_429 <= 32'h0;
    end else begin
      if (11'h1ad == _T_12323) begin
        mem_429 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_430 <= 32'h0;
    end else begin
      if (11'h1ae == _T_12323) begin
        mem_430 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_431 <= 32'h0;
    end else begin
      if (11'h1af == _T_12323) begin
        mem_431 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_432 <= 32'h0;
    end else begin
      if (11'h1b0 == _T_12323) begin
        mem_432 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_433 <= 32'h0;
    end else begin
      if (11'h1b1 == _T_12323) begin
        mem_433 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_434 <= 32'h0;
    end else begin
      if (11'h1b2 == _T_12323) begin
        mem_434 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_435 <= 32'h0;
    end else begin
      if (11'h1b3 == _T_12323) begin
        mem_435 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_436 <= 32'h0;
    end else begin
      if (11'h1b4 == _T_12323) begin
        mem_436 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_437 <= 32'h0;
    end else begin
      if (11'h1b5 == _T_12323) begin
        mem_437 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_438 <= 32'h0;
    end else begin
      if (11'h1b6 == _T_12323) begin
        mem_438 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_439 <= 32'h0;
    end else begin
      if (11'h1b7 == _T_12323) begin
        mem_439 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_440 <= 32'h0;
    end else begin
      if (11'h1b8 == _T_12323) begin
        mem_440 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_441 <= 32'h0;
    end else begin
      if (11'h1b9 == _T_12323) begin
        mem_441 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_442 <= 32'h0;
    end else begin
      if (11'h1ba == _T_12323) begin
        mem_442 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_443 <= 32'h0;
    end else begin
      if (11'h1bb == _T_12323) begin
        mem_443 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_444 <= 32'h0;
    end else begin
      if (11'h1bc == _T_12323) begin
        mem_444 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_445 <= 32'h0;
    end else begin
      if (11'h1bd == _T_12323) begin
        mem_445 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_446 <= 32'h0;
    end else begin
      if (11'h1be == _T_12323) begin
        mem_446 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_447 <= 32'h0;
    end else begin
      if (11'h1bf == _T_12323) begin
        mem_447 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_448 <= 32'h0;
    end else begin
      if (11'h1c0 == _T_12323) begin
        mem_448 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_449 <= 32'h0;
    end else begin
      if (11'h1c1 == _T_12323) begin
        mem_449 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_450 <= 32'h0;
    end else begin
      if (11'h1c2 == _T_12323) begin
        mem_450 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_451 <= 32'h0;
    end else begin
      if (11'h1c3 == _T_12323) begin
        mem_451 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_452 <= 32'h0;
    end else begin
      if (11'h1c4 == _T_12323) begin
        mem_452 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_453 <= 32'h0;
    end else begin
      if (11'h1c5 == _T_12323) begin
        mem_453 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_454 <= 32'h0;
    end else begin
      if (11'h1c6 == _T_12323) begin
        mem_454 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_455 <= 32'h0;
    end else begin
      if (11'h1c7 == _T_12323) begin
        mem_455 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_456 <= 32'h0;
    end else begin
      if (11'h1c8 == _T_12323) begin
        mem_456 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_457 <= 32'h0;
    end else begin
      if (11'h1c9 == _T_12323) begin
        mem_457 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_458 <= 32'h0;
    end else begin
      if (11'h1ca == _T_12323) begin
        mem_458 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_459 <= 32'h0;
    end else begin
      if (11'h1cb == _T_12323) begin
        mem_459 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_460 <= 32'h0;
    end else begin
      if (11'h1cc == _T_12323) begin
        mem_460 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_461 <= 32'h0;
    end else begin
      if (11'h1cd == _T_12323) begin
        mem_461 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_462 <= 32'h0;
    end else begin
      if (11'h1ce == _T_12323) begin
        mem_462 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_463 <= 32'h0;
    end else begin
      if (11'h1cf == _T_12323) begin
        mem_463 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_464 <= 32'h0;
    end else begin
      if (11'h1d0 == _T_12323) begin
        mem_464 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_465 <= 32'h0;
    end else begin
      if (11'h1d1 == _T_12323) begin
        mem_465 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_466 <= 32'h0;
    end else begin
      if (11'h1d2 == _T_12323) begin
        mem_466 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_467 <= 32'h0;
    end else begin
      if (11'h1d3 == _T_12323) begin
        mem_467 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_468 <= 32'h0;
    end else begin
      if (11'h1d4 == _T_12323) begin
        mem_468 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_469 <= 32'h0;
    end else begin
      if (11'h1d5 == _T_12323) begin
        mem_469 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_470 <= 32'h0;
    end else begin
      if (11'h1d6 == _T_12323) begin
        mem_470 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_471 <= 32'h0;
    end else begin
      if (11'h1d7 == _T_12323) begin
        mem_471 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_472 <= 32'h0;
    end else begin
      if (11'h1d8 == _T_12323) begin
        mem_472 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_473 <= 32'h0;
    end else begin
      if (11'h1d9 == _T_12323) begin
        mem_473 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_474 <= 32'h0;
    end else begin
      if (11'h1da == _T_12323) begin
        mem_474 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_475 <= 32'h0;
    end else begin
      if (11'h1db == _T_12323) begin
        mem_475 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_476 <= 32'h0;
    end else begin
      if (11'h1dc == _T_12323) begin
        mem_476 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_477 <= 32'h0;
    end else begin
      if (11'h1dd == _T_12323) begin
        mem_477 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_478 <= 32'h0;
    end else begin
      if (11'h1de == _T_12323) begin
        mem_478 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_479 <= 32'h0;
    end else begin
      if (11'h1df == _T_12323) begin
        mem_479 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_480 <= 32'h0;
    end else begin
      if (11'h1e0 == _T_12323) begin
        mem_480 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_481 <= 32'h0;
    end else begin
      if (11'h1e1 == _T_12323) begin
        mem_481 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_482 <= 32'h0;
    end else begin
      if (11'h1e2 == _T_12323) begin
        mem_482 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_483 <= 32'h0;
    end else begin
      if (11'h1e3 == _T_12323) begin
        mem_483 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_484 <= 32'h0;
    end else begin
      if (11'h1e4 == _T_12323) begin
        mem_484 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_485 <= 32'h0;
    end else begin
      if (11'h1e5 == _T_12323) begin
        mem_485 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_486 <= 32'h0;
    end else begin
      if (11'h1e6 == _T_12323) begin
        mem_486 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_487 <= 32'h0;
    end else begin
      if (11'h1e7 == _T_12323) begin
        mem_487 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_488 <= 32'h0;
    end else begin
      if (11'h1e8 == _T_12323) begin
        mem_488 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_489 <= 32'h0;
    end else begin
      if (11'h1e9 == _T_12323) begin
        mem_489 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_490 <= 32'h0;
    end else begin
      if (11'h1ea == _T_12323) begin
        mem_490 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_491 <= 32'h0;
    end else begin
      if (11'h1eb == _T_12323) begin
        mem_491 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_492 <= 32'h0;
    end else begin
      if (11'h1ec == _T_12323) begin
        mem_492 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_493 <= 32'h0;
    end else begin
      if (11'h1ed == _T_12323) begin
        mem_493 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_494 <= 32'h0;
    end else begin
      if (11'h1ee == _T_12323) begin
        mem_494 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_495 <= 32'h0;
    end else begin
      if (11'h1ef == _T_12323) begin
        mem_495 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_496 <= 32'h0;
    end else begin
      if (11'h1f0 == _T_12323) begin
        mem_496 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_497 <= 32'h0;
    end else begin
      if (11'h1f1 == _T_12323) begin
        mem_497 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_498 <= 32'h0;
    end else begin
      if (11'h1f2 == _T_12323) begin
        mem_498 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_499 <= 32'h0;
    end else begin
      if (11'h1f3 == _T_12323) begin
        mem_499 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_500 <= 32'h0;
    end else begin
      if (11'h1f4 == _T_12323) begin
        mem_500 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_501 <= 32'h0;
    end else begin
      if (11'h1f5 == _T_12323) begin
        mem_501 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_502 <= 32'h0;
    end else begin
      if (11'h1f6 == _T_12323) begin
        mem_502 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_503 <= 32'h0;
    end else begin
      if (11'h1f7 == _T_12323) begin
        mem_503 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_504 <= 32'h0;
    end else begin
      if (11'h1f8 == _T_12323) begin
        mem_504 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_505 <= 32'h0;
    end else begin
      if (11'h1f9 == _T_12323) begin
        mem_505 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_506 <= 32'h0;
    end else begin
      if (11'h1fa == _T_12323) begin
        mem_506 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_507 <= 32'h0;
    end else begin
      if (11'h1fb == _T_12323) begin
        mem_507 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_508 <= 32'h0;
    end else begin
      if (11'h1fc == _T_12323) begin
        mem_508 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_509 <= 32'h0;
    end else begin
      if (11'h1fd == _T_12323) begin
        mem_509 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_510 <= 32'h0;
    end else begin
      if (11'h1fe == _T_12323) begin
        mem_510 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_511 <= 32'h0;
    end else begin
      if (11'h1ff == _T_12323) begin
        mem_511 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_512 <= 32'h0;
    end else begin
      if (11'h200 == _T_12323) begin
        mem_512 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_513 <= 32'h0;
    end else begin
      if (11'h201 == _T_12323) begin
        mem_513 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_514 <= 32'h0;
    end else begin
      if (11'h202 == _T_12323) begin
        mem_514 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_515 <= 32'h0;
    end else begin
      if (11'h203 == _T_12323) begin
        mem_515 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_516 <= 32'h0;
    end else begin
      if (11'h204 == _T_12323) begin
        mem_516 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_517 <= 32'h0;
    end else begin
      if (11'h205 == _T_12323) begin
        mem_517 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_518 <= 32'h0;
    end else begin
      if (11'h206 == _T_12323) begin
        mem_518 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_519 <= 32'h0;
    end else begin
      if (11'h207 == _T_12323) begin
        mem_519 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_520 <= 32'h0;
    end else begin
      if (11'h208 == _T_12323) begin
        mem_520 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_521 <= 32'h0;
    end else begin
      if (11'h209 == _T_12323) begin
        mem_521 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_522 <= 32'h0;
    end else begin
      if (11'h20a == _T_12323) begin
        mem_522 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_523 <= 32'h0;
    end else begin
      if (11'h20b == _T_12323) begin
        mem_523 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_524 <= 32'h0;
    end else begin
      if (11'h20c == _T_12323) begin
        mem_524 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_525 <= 32'h0;
    end else begin
      if (11'h20d == _T_12323) begin
        mem_525 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_526 <= 32'h0;
    end else begin
      if (11'h20e == _T_12323) begin
        mem_526 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_527 <= 32'h0;
    end else begin
      if (11'h20f == _T_12323) begin
        mem_527 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_528 <= 32'h0;
    end else begin
      if (11'h210 == _T_12323) begin
        mem_528 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_529 <= 32'h0;
    end else begin
      if (11'h211 == _T_12323) begin
        mem_529 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_530 <= 32'h0;
    end else begin
      if (11'h212 == _T_12323) begin
        mem_530 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_531 <= 32'h0;
    end else begin
      if (11'h213 == _T_12323) begin
        mem_531 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_532 <= 32'h0;
    end else begin
      if (11'h214 == _T_12323) begin
        mem_532 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_533 <= 32'h0;
    end else begin
      if (11'h215 == _T_12323) begin
        mem_533 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_534 <= 32'h0;
    end else begin
      if (11'h216 == _T_12323) begin
        mem_534 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_535 <= 32'h0;
    end else begin
      if (11'h217 == _T_12323) begin
        mem_535 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_536 <= 32'h0;
    end else begin
      if (11'h218 == _T_12323) begin
        mem_536 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_537 <= 32'h0;
    end else begin
      if (11'h219 == _T_12323) begin
        mem_537 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_538 <= 32'h0;
    end else begin
      if (11'h21a == _T_12323) begin
        mem_538 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_539 <= 32'h0;
    end else begin
      if (11'h21b == _T_12323) begin
        mem_539 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_540 <= 32'h0;
    end else begin
      if (11'h21c == _T_12323) begin
        mem_540 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_541 <= 32'h0;
    end else begin
      if (11'h21d == _T_12323) begin
        mem_541 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_542 <= 32'h0;
    end else begin
      if (11'h21e == _T_12323) begin
        mem_542 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_543 <= 32'h0;
    end else begin
      if (11'h21f == _T_12323) begin
        mem_543 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_544 <= 32'h0;
    end else begin
      if (11'h220 == _T_12323) begin
        mem_544 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_545 <= 32'h0;
    end else begin
      if (11'h221 == _T_12323) begin
        mem_545 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_546 <= 32'h0;
    end else begin
      if (11'h222 == _T_12323) begin
        mem_546 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_547 <= 32'h0;
    end else begin
      if (11'h223 == _T_12323) begin
        mem_547 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_548 <= 32'h0;
    end else begin
      if (11'h224 == _T_12323) begin
        mem_548 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_549 <= 32'h0;
    end else begin
      if (11'h225 == _T_12323) begin
        mem_549 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_550 <= 32'h0;
    end else begin
      if (11'h226 == _T_12323) begin
        mem_550 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_551 <= 32'h0;
    end else begin
      if (11'h227 == _T_12323) begin
        mem_551 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_552 <= 32'h0;
    end else begin
      if (11'h228 == _T_12323) begin
        mem_552 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_553 <= 32'h0;
    end else begin
      if (11'h229 == _T_12323) begin
        mem_553 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_554 <= 32'h0;
    end else begin
      if (11'h22a == _T_12323) begin
        mem_554 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_555 <= 32'h0;
    end else begin
      if (11'h22b == _T_12323) begin
        mem_555 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_556 <= 32'h0;
    end else begin
      if (11'h22c == _T_12323) begin
        mem_556 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_557 <= 32'h0;
    end else begin
      if (11'h22d == _T_12323) begin
        mem_557 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_558 <= 32'h0;
    end else begin
      if (11'h22e == _T_12323) begin
        mem_558 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_559 <= 32'h0;
    end else begin
      if (11'h22f == _T_12323) begin
        mem_559 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_560 <= 32'h0;
    end else begin
      if (11'h230 == _T_12323) begin
        mem_560 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_561 <= 32'h0;
    end else begin
      if (11'h231 == _T_12323) begin
        mem_561 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_562 <= 32'h0;
    end else begin
      if (11'h232 == _T_12323) begin
        mem_562 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_563 <= 32'h0;
    end else begin
      if (11'h233 == _T_12323) begin
        mem_563 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_564 <= 32'h0;
    end else begin
      if (11'h234 == _T_12323) begin
        mem_564 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_565 <= 32'h0;
    end else begin
      if (11'h235 == _T_12323) begin
        mem_565 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_566 <= 32'h0;
    end else begin
      if (11'h236 == _T_12323) begin
        mem_566 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_567 <= 32'h0;
    end else begin
      if (11'h237 == _T_12323) begin
        mem_567 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_568 <= 32'h0;
    end else begin
      if (11'h238 == _T_12323) begin
        mem_568 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_569 <= 32'h0;
    end else begin
      if (11'h239 == _T_12323) begin
        mem_569 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_570 <= 32'h0;
    end else begin
      if (11'h23a == _T_12323) begin
        mem_570 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_571 <= 32'h0;
    end else begin
      if (11'h23b == _T_12323) begin
        mem_571 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_572 <= 32'h0;
    end else begin
      if (11'h23c == _T_12323) begin
        mem_572 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_573 <= 32'h0;
    end else begin
      if (11'h23d == _T_12323) begin
        mem_573 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_574 <= 32'h0;
    end else begin
      if (11'h23e == _T_12323) begin
        mem_574 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_575 <= 32'h0;
    end else begin
      if (11'h23f == _T_12323) begin
        mem_575 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_576 <= 32'h0;
    end else begin
      if (11'h240 == _T_12323) begin
        mem_576 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_577 <= 32'h0;
    end else begin
      if (11'h241 == _T_12323) begin
        mem_577 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_578 <= 32'h0;
    end else begin
      if (11'h242 == _T_12323) begin
        mem_578 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_579 <= 32'h0;
    end else begin
      if (11'h243 == _T_12323) begin
        mem_579 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_580 <= 32'h0;
    end else begin
      if (11'h244 == _T_12323) begin
        mem_580 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_581 <= 32'h0;
    end else begin
      if (11'h245 == _T_12323) begin
        mem_581 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_582 <= 32'h0;
    end else begin
      if (11'h246 == _T_12323) begin
        mem_582 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_583 <= 32'h0;
    end else begin
      if (11'h247 == _T_12323) begin
        mem_583 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_584 <= 32'h0;
    end else begin
      if (11'h248 == _T_12323) begin
        mem_584 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_585 <= 32'h0;
    end else begin
      if (11'h249 == _T_12323) begin
        mem_585 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_586 <= 32'h0;
    end else begin
      if (11'h24a == _T_12323) begin
        mem_586 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_587 <= 32'h0;
    end else begin
      if (11'h24b == _T_12323) begin
        mem_587 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_588 <= 32'h0;
    end else begin
      if (11'h24c == _T_12323) begin
        mem_588 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_589 <= 32'h0;
    end else begin
      if (11'h24d == _T_12323) begin
        mem_589 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_590 <= 32'h0;
    end else begin
      if (11'h24e == _T_12323) begin
        mem_590 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_591 <= 32'h0;
    end else begin
      if (11'h24f == _T_12323) begin
        mem_591 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_592 <= 32'h0;
    end else begin
      if (11'h250 == _T_12323) begin
        mem_592 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_593 <= 32'h0;
    end else begin
      if (11'h251 == _T_12323) begin
        mem_593 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_594 <= 32'h0;
    end else begin
      if (11'h252 == _T_12323) begin
        mem_594 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_595 <= 32'h0;
    end else begin
      if (11'h253 == _T_12323) begin
        mem_595 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_596 <= 32'h0;
    end else begin
      if (11'h254 == _T_12323) begin
        mem_596 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_597 <= 32'h0;
    end else begin
      if (11'h255 == _T_12323) begin
        mem_597 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_598 <= 32'h0;
    end else begin
      if (11'h256 == _T_12323) begin
        mem_598 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_599 <= 32'h0;
    end else begin
      if (11'h257 == _T_12323) begin
        mem_599 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_600 <= 32'h0;
    end else begin
      if (11'h258 == _T_12323) begin
        mem_600 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_601 <= 32'h0;
    end else begin
      if (11'h259 == _T_12323) begin
        mem_601 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_602 <= 32'h0;
    end else begin
      if (11'h25a == _T_12323) begin
        mem_602 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_603 <= 32'h0;
    end else begin
      if (11'h25b == _T_12323) begin
        mem_603 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_604 <= 32'h0;
    end else begin
      if (11'h25c == _T_12323) begin
        mem_604 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_605 <= 32'h0;
    end else begin
      if (11'h25d == _T_12323) begin
        mem_605 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_606 <= 32'h0;
    end else begin
      if (11'h25e == _T_12323) begin
        mem_606 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_607 <= 32'h0;
    end else begin
      if (11'h25f == _T_12323) begin
        mem_607 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_608 <= 32'h0;
    end else begin
      if (11'h260 == _T_12323) begin
        mem_608 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_609 <= 32'h0;
    end else begin
      if (11'h261 == _T_12323) begin
        mem_609 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_610 <= 32'h0;
    end else begin
      if (11'h262 == _T_12323) begin
        mem_610 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_611 <= 32'h0;
    end else begin
      if (11'h263 == _T_12323) begin
        mem_611 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_612 <= 32'h0;
    end else begin
      if (11'h264 == _T_12323) begin
        mem_612 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_613 <= 32'h0;
    end else begin
      if (11'h265 == _T_12323) begin
        mem_613 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_614 <= 32'h0;
    end else begin
      if (11'h266 == _T_12323) begin
        mem_614 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_615 <= 32'h0;
    end else begin
      if (11'h267 == _T_12323) begin
        mem_615 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_616 <= 32'h0;
    end else begin
      if (11'h268 == _T_12323) begin
        mem_616 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_617 <= 32'h0;
    end else begin
      if (11'h269 == _T_12323) begin
        mem_617 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_618 <= 32'h0;
    end else begin
      if (11'h26a == _T_12323) begin
        mem_618 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_619 <= 32'h0;
    end else begin
      if (11'h26b == _T_12323) begin
        mem_619 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_620 <= 32'h0;
    end else begin
      if (11'h26c == _T_12323) begin
        mem_620 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_621 <= 32'h0;
    end else begin
      if (11'h26d == _T_12323) begin
        mem_621 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_622 <= 32'h0;
    end else begin
      if (11'h26e == _T_12323) begin
        mem_622 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_623 <= 32'h0;
    end else begin
      if (11'h26f == _T_12323) begin
        mem_623 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_624 <= 32'h0;
    end else begin
      if (11'h270 == _T_12323) begin
        mem_624 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_625 <= 32'h0;
    end else begin
      if (11'h271 == _T_12323) begin
        mem_625 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_626 <= 32'h0;
    end else begin
      if (11'h272 == _T_12323) begin
        mem_626 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_627 <= 32'h0;
    end else begin
      if (11'h273 == _T_12323) begin
        mem_627 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_628 <= 32'h0;
    end else begin
      if (11'h274 == _T_12323) begin
        mem_628 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_629 <= 32'h0;
    end else begin
      if (11'h275 == _T_12323) begin
        mem_629 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_630 <= 32'h0;
    end else begin
      if (11'h276 == _T_12323) begin
        mem_630 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_631 <= 32'h0;
    end else begin
      if (11'h277 == _T_12323) begin
        mem_631 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_632 <= 32'h0;
    end else begin
      if (11'h278 == _T_12323) begin
        mem_632 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_633 <= 32'h0;
    end else begin
      if (11'h279 == _T_12323) begin
        mem_633 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_634 <= 32'h0;
    end else begin
      if (11'h27a == _T_12323) begin
        mem_634 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_635 <= 32'h0;
    end else begin
      if (11'h27b == _T_12323) begin
        mem_635 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_636 <= 32'h0;
    end else begin
      if (11'h27c == _T_12323) begin
        mem_636 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_637 <= 32'h0;
    end else begin
      if (11'h27d == _T_12323) begin
        mem_637 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_638 <= 32'h0;
    end else begin
      if (11'h27e == _T_12323) begin
        mem_638 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_639 <= 32'h0;
    end else begin
      if (11'h27f == _T_12323) begin
        mem_639 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_640 <= 32'h0;
    end else begin
      if (11'h280 == _T_12323) begin
        mem_640 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_641 <= 32'h0;
    end else begin
      if (11'h281 == _T_12323) begin
        mem_641 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_642 <= 32'h0;
    end else begin
      if (11'h282 == _T_12323) begin
        mem_642 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_643 <= 32'h0;
    end else begin
      if (11'h283 == _T_12323) begin
        mem_643 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_644 <= 32'h0;
    end else begin
      if (11'h284 == _T_12323) begin
        mem_644 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_645 <= 32'h0;
    end else begin
      if (11'h285 == _T_12323) begin
        mem_645 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_646 <= 32'h0;
    end else begin
      if (11'h286 == _T_12323) begin
        mem_646 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_647 <= 32'h0;
    end else begin
      if (11'h287 == _T_12323) begin
        mem_647 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_648 <= 32'h0;
    end else begin
      if (11'h288 == _T_12323) begin
        mem_648 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_649 <= 32'h0;
    end else begin
      if (11'h289 == _T_12323) begin
        mem_649 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_650 <= 32'h0;
    end else begin
      if (11'h28a == _T_12323) begin
        mem_650 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_651 <= 32'h0;
    end else begin
      if (11'h28b == _T_12323) begin
        mem_651 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_652 <= 32'h0;
    end else begin
      if (11'h28c == _T_12323) begin
        mem_652 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_653 <= 32'h0;
    end else begin
      if (11'h28d == _T_12323) begin
        mem_653 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_654 <= 32'h0;
    end else begin
      if (11'h28e == _T_12323) begin
        mem_654 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_655 <= 32'h0;
    end else begin
      if (11'h28f == _T_12323) begin
        mem_655 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_656 <= 32'h0;
    end else begin
      if (11'h290 == _T_12323) begin
        mem_656 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_657 <= 32'h0;
    end else begin
      if (11'h291 == _T_12323) begin
        mem_657 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_658 <= 32'h0;
    end else begin
      if (11'h292 == _T_12323) begin
        mem_658 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_659 <= 32'h0;
    end else begin
      if (11'h293 == _T_12323) begin
        mem_659 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_660 <= 32'h0;
    end else begin
      if (11'h294 == _T_12323) begin
        mem_660 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_661 <= 32'h0;
    end else begin
      if (11'h295 == _T_12323) begin
        mem_661 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_662 <= 32'h0;
    end else begin
      if (11'h296 == _T_12323) begin
        mem_662 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_663 <= 32'h0;
    end else begin
      if (11'h297 == _T_12323) begin
        mem_663 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_664 <= 32'h0;
    end else begin
      if (11'h298 == _T_12323) begin
        mem_664 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_665 <= 32'h0;
    end else begin
      if (11'h299 == _T_12323) begin
        mem_665 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_666 <= 32'h0;
    end else begin
      if (11'h29a == _T_12323) begin
        mem_666 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_667 <= 32'h0;
    end else begin
      if (11'h29b == _T_12323) begin
        mem_667 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_668 <= 32'h0;
    end else begin
      if (11'h29c == _T_12323) begin
        mem_668 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_669 <= 32'h0;
    end else begin
      if (11'h29d == _T_12323) begin
        mem_669 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_670 <= 32'h0;
    end else begin
      if (11'h29e == _T_12323) begin
        mem_670 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_671 <= 32'h0;
    end else begin
      if (11'h29f == _T_12323) begin
        mem_671 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_672 <= 32'h0;
    end else begin
      if (11'h2a0 == _T_12323) begin
        mem_672 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_673 <= 32'h0;
    end else begin
      if (11'h2a1 == _T_12323) begin
        mem_673 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_674 <= 32'h0;
    end else begin
      if (11'h2a2 == _T_12323) begin
        mem_674 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_675 <= 32'h0;
    end else begin
      if (11'h2a3 == _T_12323) begin
        mem_675 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_676 <= 32'h0;
    end else begin
      if (11'h2a4 == _T_12323) begin
        mem_676 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_677 <= 32'h0;
    end else begin
      if (11'h2a5 == _T_12323) begin
        mem_677 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_678 <= 32'h0;
    end else begin
      if (11'h2a6 == _T_12323) begin
        mem_678 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_679 <= 32'h0;
    end else begin
      if (11'h2a7 == _T_12323) begin
        mem_679 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_680 <= 32'h0;
    end else begin
      if (11'h2a8 == _T_12323) begin
        mem_680 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_681 <= 32'h0;
    end else begin
      if (11'h2a9 == _T_12323) begin
        mem_681 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_682 <= 32'h0;
    end else begin
      if (11'h2aa == _T_12323) begin
        mem_682 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_683 <= 32'h0;
    end else begin
      if (11'h2ab == _T_12323) begin
        mem_683 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_684 <= 32'h0;
    end else begin
      if (11'h2ac == _T_12323) begin
        mem_684 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_685 <= 32'h0;
    end else begin
      if (11'h2ad == _T_12323) begin
        mem_685 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_686 <= 32'h0;
    end else begin
      if (11'h2ae == _T_12323) begin
        mem_686 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_687 <= 32'h0;
    end else begin
      if (11'h2af == _T_12323) begin
        mem_687 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_688 <= 32'h0;
    end else begin
      if (11'h2b0 == _T_12323) begin
        mem_688 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_689 <= 32'h0;
    end else begin
      if (11'h2b1 == _T_12323) begin
        mem_689 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_690 <= 32'h0;
    end else begin
      if (11'h2b2 == _T_12323) begin
        mem_690 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_691 <= 32'h0;
    end else begin
      if (11'h2b3 == _T_12323) begin
        mem_691 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_692 <= 32'h0;
    end else begin
      if (11'h2b4 == _T_12323) begin
        mem_692 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_693 <= 32'h0;
    end else begin
      if (11'h2b5 == _T_12323) begin
        mem_693 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_694 <= 32'h0;
    end else begin
      if (11'h2b6 == _T_12323) begin
        mem_694 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_695 <= 32'h0;
    end else begin
      if (11'h2b7 == _T_12323) begin
        mem_695 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_696 <= 32'h0;
    end else begin
      if (11'h2b8 == _T_12323) begin
        mem_696 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_697 <= 32'h0;
    end else begin
      if (11'h2b9 == _T_12323) begin
        mem_697 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_698 <= 32'h0;
    end else begin
      if (11'h2ba == _T_12323) begin
        mem_698 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_699 <= 32'h0;
    end else begin
      if (11'h2bb == _T_12323) begin
        mem_699 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_700 <= 32'h0;
    end else begin
      if (11'h2bc == _T_12323) begin
        mem_700 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_701 <= 32'h0;
    end else begin
      if (11'h2bd == _T_12323) begin
        mem_701 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_702 <= 32'h0;
    end else begin
      if (11'h2be == _T_12323) begin
        mem_702 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_703 <= 32'h0;
    end else begin
      if (11'h2bf == _T_12323) begin
        mem_703 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_704 <= 32'h0;
    end else begin
      if (11'h2c0 == _T_12323) begin
        mem_704 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_705 <= 32'h0;
    end else begin
      if (11'h2c1 == _T_12323) begin
        mem_705 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_706 <= 32'h0;
    end else begin
      if (11'h2c2 == _T_12323) begin
        mem_706 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_707 <= 32'h0;
    end else begin
      if (11'h2c3 == _T_12323) begin
        mem_707 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_708 <= 32'h0;
    end else begin
      if (11'h2c4 == _T_12323) begin
        mem_708 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_709 <= 32'h0;
    end else begin
      if (11'h2c5 == _T_12323) begin
        mem_709 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_710 <= 32'h0;
    end else begin
      if (11'h2c6 == _T_12323) begin
        mem_710 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_711 <= 32'h0;
    end else begin
      if (11'h2c7 == _T_12323) begin
        mem_711 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_712 <= 32'h0;
    end else begin
      if (11'h2c8 == _T_12323) begin
        mem_712 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_713 <= 32'h0;
    end else begin
      if (11'h2c9 == _T_12323) begin
        mem_713 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_714 <= 32'h0;
    end else begin
      if (11'h2ca == _T_12323) begin
        mem_714 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_715 <= 32'h0;
    end else begin
      if (11'h2cb == _T_12323) begin
        mem_715 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_716 <= 32'h0;
    end else begin
      if (11'h2cc == _T_12323) begin
        mem_716 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_717 <= 32'h0;
    end else begin
      if (11'h2cd == _T_12323) begin
        mem_717 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_718 <= 32'h0;
    end else begin
      if (11'h2ce == _T_12323) begin
        mem_718 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_719 <= 32'h0;
    end else begin
      if (11'h2cf == _T_12323) begin
        mem_719 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_720 <= 32'h0;
    end else begin
      if (11'h2d0 == _T_12323) begin
        mem_720 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_721 <= 32'h0;
    end else begin
      if (11'h2d1 == _T_12323) begin
        mem_721 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_722 <= 32'h0;
    end else begin
      if (11'h2d2 == _T_12323) begin
        mem_722 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_723 <= 32'h0;
    end else begin
      if (11'h2d3 == _T_12323) begin
        mem_723 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_724 <= 32'h0;
    end else begin
      if (11'h2d4 == _T_12323) begin
        mem_724 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_725 <= 32'h0;
    end else begin
      if (11'h2d5 == _T_12323) begin
        mem_725 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_726 <= 32'h0;
    end else begin
      if (11'h2d6 == _T_12323) begin
        mem_726 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_727 <= 32'h0;
    end else begin
      if (11'h2d7 == _T_12323) begin
        mem_727 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_728 <= 32'h0;
    end else begin
      if (11'h2d8 == _T_12323) begin
        mem_728 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_729 <= 32'h0;
    end else begin
      if (11'h2d9 == _T_12323) begin
        mem_729 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_730 <= 32'h0;
    end else begin
      if (11'h2da == _T_12323) begin
        mem_730 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_731 <= 32'h0;
    end else begin
      if (11'h2db == _T_12323) begin
        mem_731 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_732 <= 32'h0;
    end else begin
      if (11'h2dc == _T_12323) begin
        mem_732 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_733 <= 32'h0;
    end else begin
      if (11'h2dd == _T_12323) begin
        mem_733 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_734 <= 32'h0;
    end else begin
      if (11'h2de == _T_12323) begin
        mem_734 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_735 <= 32'h0;
    end else begin
      if (11'h2df == _T_12323) begin
        mem_735 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_736 <= 32'h0;
    end else begin
      if (11'h2e0 == _T_12323) begin
        mem_736 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_737 <= 32'h0;
    end else begin
      if (11'h2e1 == _T_12323) begin
        mem_737 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_738 <= 32'h0;
    end else begin
      if (11'h2e2 == _T_12323) begin
        mem_738 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_739 <= 32'h0;
    end else begin
      if (11'h2e3 == _T_12323) begin
        mem_739 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_740 <= 32'h0;
    end else begin
      if (11'h2e4 == _T_12323) begin
        mem_740 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_741 <= 32'h0;
    end else begin
      if (11'h2e5 == _T_12323) begin
        mem_741 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_742 <= 32'h0;
    end else begin
      if (11'h2e6 == _T_12323) begin
        mem_742 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_743 <= 32'h0;
    end else begin
      if (11'h2e7 == _T_12323) begin
        mem_743 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_744 <= 32'h0;
    end else begin
      if (11'h2e8 == _T_12323) begin
        mem_744 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_745 <= 32'h0;
    end else begin
      if (11'h2e9 == _T_12323) begin
        mem_745 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_746 <= 32'h0;
    end else begin
      if (11'h2ea == _T_12323) begin
        mem_746 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_747 <= 32'h0;
    end else begin
      if (11'h2eb == _T_12323) begin
        mem_747 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_748 <= 32'h0;
    end else begin
      if (11'h2ec == _T_12323) begin
        mem_748 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_749 <= 32'h0;
    end else begin
      if (11'h2ed == _T_12323) begin
        mem_749 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_750 <= 32'h0;
    end else begin
      if (11'h2ee == _T_12323) begin
        mem_750 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_751 <= 32'h0;
    end else begin
      if (11'h2ef == _T_12323) begin
        mem_751 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_752 <= 32'h0;
    end else begin
      if (11'h2f0 == _T_12323) begin
        mem_752 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_753 <= 32'h0;
    end else begin
      if (11'h2f1 == _T_12323) begin
        mem_753 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_754 <= 32'h0;
    end else begin
      if (11'h2f2 == _T_12323) begin
        mem_754 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_755 <= 32'h0;
    end else begin
      if (11'h2f3 == _T_12323) begin
        mem_755 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_756 <= 32'h0;
    end else begin
      if (11'h2f4 == _T_12323) begin
        mem_756 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_757 <= 32'h0;
    end else begin
      if (11'h2f5 == _T_12323) begin
        mem_757 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_758 <= 32'h0;
    end else begin
      if (11'h2f6 == _T_12323) begin
        mem_758 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_759 <= 32'h0;
    end else begin
      if (11'h2f7 == _T_12323) begin
        mem_759 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_760 <= 32'h0;
    end else begin
      if (11'h2f8 == _T_12323) begin
        mem_760 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_761 <= 32'h0;
    end else begin
      if (11'h2f9 == _T_12323) begin
        mem_761 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_762 <= 32'h0;
    end else begin
      if (11'h2fa == _T_12323) begin
        mem_762 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_763 <= 32'h0;
    end else begin
      if (11'h2fb == _T_12323) begin
        mem_763 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_764 <= 32'h0;
    end else begin
      if (11'h2fc == _T_12323) begin
        mem_764 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_765 <= 32'h0;
    end else begin
      if (11'h2fd == _T_12323) begin
        mem_765 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_766 <= 32'h0;
    end else begin
      if (11'h2fe == _T_12323) begin
        mem_766 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_767 <= 32'h0;
    end else begin
      if (11'h2ff == _T_12323) begin
        mem_767 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_768 <= 32'h0;
    end else begin
      if (11'h300 == _T_12323) begin
        mem_768 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_769 <= 32'h0;
    end else begin
      if (11'h301 == _T_12323) begin
        mem_769 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_770 <= 32'h0;
    end else begin
      if (11'h302 == _T_12323) begin
        mem_770 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_771 <= 32'h0;
    end else begin
      if (11'h303 == _T_12323) begin
        mem_771 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_772 <= 32'h0;
    end else begin
      if (11'h304 == _T_12323) begin
        mem_772 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_773 <= 32'h0;
    end else begin
      if (11'h305 == _T_12323) begin
        mem_773 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_774 <= 32'h0;
    end else begin
      if (11'h306 == _T_12323) begin
        mem_774 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_775 <= 32'h0;
    end else begin
      if (11'h307 == _T_12323) begin
        mem_775 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_776 <= 32'h0;
    end else begin
      if (11'h308 == _T_12323) begin
        mem_776 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_777 <= 32'h0;
    end else begin
      if (11'h309 == _T_12323) begin
        mem_777 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_778 <= 32'h0;
    end else begin
      if (11'h30a == _T_12323) begin
        mem_778 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_779 <= 32'h0;
    end else begin
      if (11'h30b == _T_12323) begin
        mem_779 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_780 <= 32'h0;
    end else begin
      if (11'h30c == _T_12323) begin
        mem_780 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_781 <= 32'h0;
    end else begin
      if (11'h30d == _T_12323) begin
        mem_781 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_782 <= 32'h0;
    end else begin
      if (11'h30e == _T_12323) begin
        mem_782 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_783 <= 32'h0;
    end else begin
      if (11'h30f == _T_12323) begin
        mem_783 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_784 <= 32'h0;
    end else begin
      if (11'h310 == _T_12323) begin
        mem_784 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_785 <= 32'h0;
    end else begin
      if (11'h311 == _T_12323) begin
        mem_785 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_786 <= 32'h0;
    end else begin
      if (11'h312 == _T_12323) begin
        mem_786 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_787 <= 32'h0;
    end else begin
      if (11'h313 == _T_12323) begin
        mem_787 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_788 <= 32'h0;
    end else begin
      if (11'h314 == _T_12323) begin
        mem_788 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_789 <= 32'h0;
    end else begin
      if (11'h315 == _T_12323) begin
        mem_789 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_790 <= 32'h0;
    end else begin
      if (11'h316 == _T_12323) begin
        mem_790 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_791 <= 32'h0;
    end else begin
      if (11'h317 == _T_12323) begin
        mem_791 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_792 <= 32'h0;
    end else begin
      if (11'h318 == _T_12323) begin
        mem_792 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_793 <= 32'h0;
    end else begin
      if (11'h319 == _T_12323) begin
        mem_793 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_794 <= 32'h0;
    end else begin
      if (11'h31a == _T_12323) begin
        mem_794 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_795 <= 32'h0;
    end else begin
      if (11'h31b == _T_12323) begin
        mem_795 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_796 <= 32'h0;
    end else begin
      if (11'h31c == _T_12323) begin
        mem_796 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_797 <= 32'h0;
    end else begin
      if (11'h31d == _T_12323) begin
        mem_797 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_798 <= 32'h0;
    end else begin
      if (11'h31e == _T_12323) begin
        mem_798 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_799 <= 32'h0;
    end else begin
      if (11'h31f == _T_12323) begin
        mem_799 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_800 <= 32'h0;
    end else begin
      if (11'h320 == _T_12323) begin
        mem_800 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_801 <= 32'h0;
    end else begin
      if (11'h321 == _T_12323) begin
        mem_801 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_802 <= 32'h0;
    end else begin
      if (11'h322 == _T_12323) begin
        mem_802 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_803 <= 32'h0;
    end else begin
      if (11'h323 == _T_12323) begin
        mem_803 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_804 <= 32'h0;
    end else begin
      if (11'h324 == _T_12323) begin
        mem_804 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_805 <= 32'h0;
    end else begin
      if (11'h325 == _T_12323) begin
        mem_805 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_806 <= 32'h0;
    end else begin
      if (11'h326 == _T_12323) begin
        mem_806 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_807 <= 32'h0;
    end else begin
      if (11'h327 == _T_12323) begin
        mem_807 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_808 <= 32'h0;
    end else begin
      if (11'h328 == _T_12323) begin
        mem_808 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_809 <= 32'h0;
    end else begin
      if (11'h329 == _T_12323) begin
        mem_809 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_810 <= 32'h0;
    end else begin
      if (11'h32a == _T_12323) begin
        mem_810 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_811 <= 32'h0;
    end else begin
      if (11'h32b == _T_12323) begin
        mem_811 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_812 <= 32'h0;
    end else begin
      if (11'h32c == _T_12323) begin
        mem_812 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_813 <= 32'h0;
    end else begin
      if (11'h32d == _T_12323) begin
        mem_813 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_814 <= 32'h0;
    end else begin
      if (11'h32e == _T_12323) begin
        mem_814 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_815 <= 32'h0;
    end else begin
      if (11'h32f == _T_12323) begin
        mem_815 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_816 <= 32'h0;
    end else begin
      if (11'h330 == _T_12323) begin
        mem_816 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_817 <= 32'h0;
    end else begin
      if (11'h331 == _T_12323) begin
        mem_817 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_818 <= 32'h0;
    end else begin
      if (11'h332 == _T_12323) begin
        mem_818 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_819 <= 32'h0;
    end else begin
      if (11'h333 == _T_12323) begin
        mem_819 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_820 <= 32'h0;
    end else begin
      if (11'h334 == _T_12323) begin
        mem_820 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_821 <= 32'h0;
    end else begin
      if (11'h335 == _T_12323) begin
        mem_821 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_822 <= 32'h0;
    end else begin
      if (11'h336 == _T_12323) begin
        mem_822 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_823 <= 32'h0;
    end else begin
      if (11'h337 == _T_12323) begin
        mem_823 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_824 <= 32'h0;
    end else begin
      if (11'h338 == _T_12323) begin
        mem_824 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_825 <= 32'h0;
    end else begin
      if (11'h339 == _T_12323) begin
        mem_825 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_826 <= 32'h0;
    end else begin
      if (11'h33a == _T_12323) begin
        mem_826 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_827 <= 32'h0;
    end else begin
      if (11'h33b == _T_12323) begin
        mem_827 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_828 <= 32'h0;
    end else begin
      if (11'h33c == _T_12323) begin
        mem_828 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_829 <= 32'h0;
    end else begin
      if (11'h33d == _T_12323) begin
        mem_829 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_830 <= 32'h0;
    end else begin
      if (11'h33e == _T_12323) begin
        mem_830 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_831 <= 32'h0;
    end else begin
      if (11'h33f == _T_12323) begin
        mem_831 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_832 <= 32'h0;
    end else begin
      if (11'h340 == _T_12323) begin
        mem_832 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_833 <= 32'h0;
    end else begin
      if (11'h341 == _T_12323) begin
        mem_833 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_834 <= 32'h0;
    end else begin
      if (11'h342 == _T_12323) begin
        mem_834 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_835 <= 32'h0;
    end else begin
      if (11'h343 == _T_12323) begin
        mem_835 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_836 <= 32'h0;
    end else begin
      if (11'h344 == _T_12323) begin
        mem_836 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_837 <= 32'h0;
    end else begin
      if (11'h345 == _T_12323) begin
        mem_837 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_838 <= 32'h0;
    end else begin
      if (11'h346 == _T_12323) begin
        mem_838 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_839 <= 32'h0;
    end else begin
      if (11'h347 == _T_12323) begin
        mem_839 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_840 <= 32'h0;
    end else begin
      if (11'h348 == _T_12323) begin
        mem_840 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_841 <= 32'h0;
    end else begin
      if (11'h349 == _T_12323) begin
        mem_841 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_842 <= 32'h0;
    end else begin
      if (11'h34a == _T_12323) begin
        mem_842 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_843 <= 32'h0;
    end else begin
      if (11'h34b == _T_12323) begin
        mem_843 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_844 <= 32'h0;
    end else begin
      if (11'h34c == _T_12323) begin
        mem_844 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_845 <= 32'h0;
    end else begin
      if (11'h34d == _T_12323) begin
        mem_845 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_846 <= 32'h0;
    end else begin
      if (11'h34e == _T_12323) begin
        mem_846 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_847 <= 32'h0;
    end else begin
      if (11'h34f == _T_12323) begin
        mem_847 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_848 <= 32'h0;
    end else begin
      if (11'h350 == _T_12323) begin
        mem_848 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_849 <= 32'h0;
    end else begin
      if (11'h351 == _T_12323) begin
        mem_849 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_850 <= 32'h0;
    end else begin
      if (11'h352 == _T_12323) begin
        mem_850 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_851 <= 32'h0;
    end else begin
      if (11'h353 == _T_12323) begin
        mem_851 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_852 <= 32'h0;
    end else begin
      if (11'h354 == _T_12323) begin
        mem_852 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_853 <= 32'h0;
    end else begin
      if (11'h355 == _T_12323) begin
        mem_853 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_854 <= 32'h0;
    end else begin
      if (11'h356 == _T_12323) begin
        mem_854 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_855 <= 32'h0;
    end else begin
      if (11'h357 == _T_12323) begin
        mem_855 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_856 <= 32'h0;
    end else begin
      if (11'h358 == _T_12323) begin
        mem_856 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_857 <= 32'h0;
    end else begin
      if (11'h359 == _T_12323) begin
        mem_857 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_858 <= 32'h0;
    end else begin
      if (11'h35a == _T_12323) begin
        mem_858 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_859 <= 32'h0;
    end else begin
      if (11'h35b == _T_12323) begin
        mem_859 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_860 <= 32'h0;
    end else begin
      if (11'h35c == _T_12323) begin
        mem_860 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_861 <= 32'h0;
    end else begin
      if (11'h35d == _T_12323) begin
        mem_861 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_862 <= 32'h0;
    end else begin
      if (11'h35e == _T_12323) begin
        mem_862 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_863 <= 32'h0;
    end else begin
      if (11'h35f == _T_12323) begin
        mem_863 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_864 <= 32'h0;
    end else begin
      if (11'h360 == _T_12323) begin
        mem_864 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_865 <= 32'h0;
    end else begin
      if (11'h361 == _T_12323) begin
        mem_865 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_866 <= 32'h0;
    end else begin
      if (11'h362 == _T_12323) begin
        mem_866 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_867 <= 32'h0;
    end else begin
      if (11'h363 == _T_12323) begin
        mem_867 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_868 <= 32'h0;
    end else begin
      if (11'h364 == _T_12323) begin
        mem_868 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_869 <= 32'h0;
    end else begin
      if (11'h365 == _T_12323) begin
        mem_869 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_870 <= 32'h0;
    end else begin
      if (11'h366 == _T_12323) begin
        mem_870 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_871 <= 32'h0;
    end else begin
      if (11'h367 == _T_12323) begin
        mem_871 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_872 <= 32'h0;
    end else begin
      if (11'h368 == _T_12323) begin
        mem_872 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_873 <= 32'h0;
    end else begin
      if (11'h369 == _T_12323) begin
        mem_873 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_874 <= 32'h0;
    end else begin
      if (11'h36a == _T_12323) begin
        mem_874 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_875 <= 32'h0;
    end else begin
      if (11'h36b == _T_12323) begin
        mem_875 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_876 <= 32'h0;
    end else begin
      if (11'h36c == _T_12323) begin
        mem_876 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_877 <= 32'h0;
    end else begin
      if (11'h36d == _T_12323) begin
        mem_877 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_878 <= 32'h0;
    end else begin
      if (11'h36e == _T_12323) begin
        mem_878 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_879 <= 32'h0;
    end else begin
      if (11'h36f == _T_12323) begin
        mem_879 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_880 <= 32'h0;
    end else begin
      if (11'h370 == _T_12323) begin
        mem_880 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_881 <= 32'h0;
    end else begin
      if (11'h371 == _T_12323) begin
        mem_881 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_882 <= 32'h0;
    end else begin
      if (11'h372 == _T_12323) begin
        mem_882 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_883 <= 32'h0;
    end else begin
      if (11'h373 == _T_12323) begin
        mem_883 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_884 <= 32'h0;
    end else begin
      if (11'h374 == _T_12323) begin
        mem_884 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_885 <= 32'h0;
    end else begin
      if (11'h375 == _T_12323) begin
        mem_885 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_886 <= 32'h0;
    end else begin
      if (11'h376 == _T_12323) begin
        mem_886 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_887 <= 32'h0;
    end else begin
      if (11'h377 == _T_12323) begin
        mem_887 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_888 <= 32'h0;
    end else begin
      if (11'h378 == _T_12323) begin
        mem_888 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_889 <= 32'h0;
    end else begin
      if (11'h379 == _T_12323) begin
        mem_889 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_890 <= 32'h0;
    end else begin
      if (11'h37a == _T_12323) begin
        mem_890 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_891 <= 32'h0;
    end else begin
      if (11'h37b == _T_12323) begin
        mem_891 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_892 <= 32'h0;
    end else begin
      if (11'h37c == _T_12323) begin
        mem_892 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_893 <= 32'h0;
    end else begin
      if (11'h37d == _T_12323) begin
        mem_893 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_894 <= 32'h0;
    end else begin
      if (11'h37e == _T_12323) begin
        mem_894 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_895 <= 32'h0;
    end else begin
      if (11'h37f == _T_12323) begin
        mem_895 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_896 <= 32'h0;
    end else begin
      if (11'h380 == _T_12323) begin
        mem_896 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_897 <= 32'h0;
    end else begin
      if (11'h381 == _T_12323) begin
        mem_897 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_898 <= 32'h0;
    end else begin
      if (11'h382 == _T_12323) begin
        mem_898 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_899 <= 32'h0;
    end else begin
      if (11'h383 == _T_12323) begin
        mem_899 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_900 <= 32'h0;
    end else begin
      if (11'h384 == _T_12323) begin
        mem_900 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_901 <= 32'h0;
    end else begin
      if (11'h385 == _T_12323) begin
        mem_901 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_902 <= 32'h0;
    end else begin
      if (11'h386 == _T_12323) begin
        mem_902 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_903 <= 32'h0;
    end else begin
      if (11'h387 == _T_12323) begin
        mem_903 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_904 <= 32'h0;
    end else begin
      if (11'h388 == _T_12323) begin
        mem_904 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_905 <= 32'h0;
    end else begin
      if (11'h389 == _T_12323) begin
        mem_905 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_906 <= 32'h0;
    end else begin
      if (11'h38a == _T_12323) begin
        mem_906 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_907 <= 32'h0;
    end else begin
      if (11'h38b == _T_12323) begin
        mem_907 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_908 <= 32'h0;
    end else begin
      if (11'h38c == _T_12323) begin
        mem_908 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_909 <= 32'h0;
    end else begin
      if (11'h38d == _T_12323) begin
        mem_909 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_910 <= 32'h0;
    end else begin
      if (11'h38e == _T_12323) begin
        mem_910 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_911 <= 32'h0;
    end else begin
      if (11'h38f == _T_12323) begin
        mem_911 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_912 <= 32'h0;
    end else begin
      if (11'h390 == _T_12323) begin
        mem_912 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_913 <= 32'h0;
    end else begin
      if (11'h391 == _T_12323) begin
        mem_913 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_914 <= 32'h0;
    end else begin
      if (11'h392 == _T_12323) begin
        mem_914 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_915 <= 32'h0;
    end else begin
      if (11'h393 == _T_12323) begin
        mem_915 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_916 <= 32'h0;
    end else begin
      if (11'h394 == _T_12323) begin
        mem_916 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_917 <= 32'h0;
    end else begin
      if (11'h395 == _T_12323) begin
        mem_917 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_918 <= 32'h0;
    end else begin
      if (11'h396 == _T_12323) begin
        mem_918 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_919 <= 32'h0;
    end else begin
      if (11'h397 == _T_12323) begin
        mem_919 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_920 <= 32'h0;
    end else begin
      if (11'h398 == _T_12323) begin
        mem_920 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_921 <= 32'h0;
    end else begin
      if (11'h399 == _T_12323) begin
        mem_921 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_922 <= 32'h0;
    end else begin
      if (11'h39a == _T_12323) begin
        mem_922 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_923 <= 32'h0;
    end else begin
      if (11'h39b == _T_12323) begin
        mem_923 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_924 <= 32'h0;
    end else begin
      if (11'h39c == _T_12323) begin
        mem_924 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_925 <= 32'h0;
    end else begin
      if (11'h39d == _T_12323) begin
        mem_925 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_926 <= 32'h0;
    end else begin
      if (11'h39e == _T_12323) begin
        mem_926 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_927 <= 32'h0;
    end else begin
      if (11'h39f == _T_12323) begin
        mem_927 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_928 <= 32'h0;
    end else begin
      if (11'h3a0 == _T_12323) begin
        mem_928 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_929 <= 32'h0;
    end else begin
      if (11'h3a1 == _T_12323) begin
        mem_929 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_930 <= 32'h0;
    end else begin
      if (11'h3a2 == _T_12323) begin
        mem_930 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_931 <= 32'h0;
    end else begin
      if (11'h3a3 == _T_12323) begin
        mem_931 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_932 <= 32'h0;
    end else begin
      if (11'h3a4 == _T_12323) begin
        mem_932 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_933 <= 32'h0;
    end else begin
      if (11'h3a5 == _T_12323) begin
        mem_933 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_934 <= 32'h0;
    end else begin
      if (11'h3a6 == _T_12323) begin
        mem_934 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_935 <= 32'h0;
    end else begin
      if (11'h3a7 == _T_12323) begin
        mem_935 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_936 <= 32'h0;
    end else begin
      if (11'h3a8 == _T_12323) begin
        mem_936 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_937 <= 32'h0;
    end else begin
      if (11'h3a9 == _T_12323) begin
        mem_937 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_938 <= 32'h0;
    end else begin
      if (11'h3aa == _T_12323) begin
        mem_938 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_939 <= 32'h0;
    end else begin
      if (11'h3ab == _T_12323) begin
        mem_939 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_940 <= 32'h0;
    end else begin
      if (11'h3ac == _T_12323) begin
        mem_940 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_941 <= 32'h0;
    end else begin
      if (11'h3ad == _T_12323) begin
        mem_941 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_942 <= 32'h0;
    end else begin
      if (11'h3ae == _T_12323) begin
        mem_942 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_943 <= 32'h0;
    end else begin
      if (11'h3af == _T_12323) begin
        mem_943 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_944 <= 32'h0;
    end else begin
      if (11'h3b0 == _T_12323) begin
        mem_944 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_945 <= 32'h0;
    end else begin
      if (11'h3b1 == _T_12323) begin
        mem_945 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_946 <= 32'h0;
    end else begin
      if (11'h3b2 == _T_12323) begin
        mem_946 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_947 <= 32'h0;
    end else begin
      if (11'h3b3 == _T_12323) begin
        mem_947 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_948 <= 32'h0;
    end else begin
      if (11'h3b4 == _T_12323) begin
        mem_948 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_949 <= 32'h0;
    end else begin
      if (11'h3b5 == _T_12323) begin
        mem_949 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_950 <= 32'h0;
    end else begin
      if (11'h3b6 == _T_12323) begin
        mem_950 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_951 <= 32'h0;
    end else begin
      if (11'h3b7 == _T_12323) begin
        mem_951 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_952 <= 32'h0;
    end else begin
      if (11'h3b8 == _T_12323) begin
        mem_952 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_953 <= 32'h0;
    end else begin
      if (11'h3b9 == _T_12323) begin
        mem_953 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_954 <= 32'h0;
    end else begin
      if (11'h3ba == _T_12323) begin
        mem_954 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_955 <= 32'h0;
    end else begin
      if (11'h3bb == _T_12323) begin
        mem_955 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_956 <= 32'h0;
    end else begin
      if (11'h3bc == _T_12323) begin
        mem_956 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_957 <= 32'h0;
    end else begin
      if (11'h3bd == _T_12323) begin
        mem_957 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_958 <= 32'h0;
    end else begin
      if (11'h3be == _T_12323) begin
        mem_958 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_959 <= 32'h0;
    end else begin
      if (11'h3bf == _T_12323) begin
        mem_959 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_960 <= 32'h0;
    end else begin
      if (11'h3c0 == _T_12323) begin
        mem_960 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_961 <= 32'h0;
    end else begin
      if (11'h3c1 == _T_12323) begin
        mem_961 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_962 <= 32'h0;
    end else begin
      if (11'h3c2 == _T_12323) begin
        mem_962 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_963 <= 32'h0;
    end else begin
      if (11'h3c3 == _T_12323) begin
        mem_963 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_964 <= 32'h0;
    end else begin
      if (11'h3c4 == _T_12323) begin
        mem_964 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_965 <= 32'h0;
    end else begin
      if (11'h3c5 == _T_12323) begin
        mem_965 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_966 <= 32'h0;
    end else begin
      if (11'h3c6 == _T_12323) begin
        mem_966 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_967 <= 32'h0;
    end else begin
      if (11'h3c7 == _T_12323) begin
        mem_967 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_968 <= 32'h0;
    end else begin
      if (11'h3c8 == _T_12323) begin
        mem_968 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_969 <= 32'h0;
    end else begin
      if (11'h3c9 == _T_12323) begin
        mem_969 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_970 <= 32'h0;
    end else begin
      if (11'h3ca == _T_12323) begin
        mem_970 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_971 <= 32'h0;
    end else begin
      if (11'h3cb == _T_12323) begin
        mem_971 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_972 <= 32'h0;
    end else begin
      if (11'h3cc == _T_12323) begin
        mem_972 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_973 <= 32'h0;
    end else begin
      if (11'h3cd == _T_12323) begin
        mem_973 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_974 <= 32'h0;
    end else begin
      if (11'h3ce == _T_12323) begin
        mem_974 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_975 <= 32'h0;
    end else begin
      if (11'h3cf == _T_12323) begin
        mem_975 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_976 <= 32'h0;
    end else begin
      if (11'h3d0 == _T_12323) begin
        mem_976 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_977 <= 32'h0;
    end else begin
      if (11'h3d1 == _T_12323) begin
        mem_977 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_978 <= 32'h0;
    end else begin
      if (11'h3d2 == _T_12323) begin
        mem_978 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_979 <= 32'h0;
    end else begin
      if (11'h3d3 == _T_12323) begin
        mem_979 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_980 <= 32'h0;
    end else begin
      if (11'h3d4 == _T_12323) begin
        mem_980 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_981 <= 32'h0;
    end else begin
      if (11'h3d5 == _T_12323) begin
        mem_981 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_982 <= 32'h0;
    end else begin
      if (11'h3d6 == _T_12323) begin
        mem_982 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_983 <= 32'h0;
    end else begin
      if (11'h3d7 == _T_12323) begin
        mem_983 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_984 <= 32'h0;
    end else begin
      if (11'h3d8 == _T_12323) begin
        mem_984 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_985 <= 32'h0;
    end else begin
      if (11'h3d9 == _T_12323) begin
        mem_985 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_986 <= 32'h0;
    end else begin
      if (11'h3da == _T_12323) begin
        mem_986 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_987 <= 32'h0;
    end else begin
      if (11'h3db == _T_12323) begin
        mem_987 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_988 <= 32'h0;
    end else begin
      if (11'h3dc == _T_12323) begin
        mem_988 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_989 <= 32'h0;
    end else begin
      if (11'h3dd == _T_12323) begin
        mem_989 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_990 <= 32'h0;
    end else begin
      if (11'h3de == _T_12323) begin
        mem_990 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_991 <= 32'h0;
    end else begin
      if (11'h3df == _T_12323) begin
        mem_991 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_992 <= 32'h0;
    end else begin
      if (11'h3e0 == _T_12323) begin
        mem_992 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_993 <= 32'h0;
    end else begin
      if (11'h3e1 == _T_12323) begin
        mem_993 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_994 <= 32'h0;
    end else begin
      if (11'h3e2 == _T_12323) begin
        mem_994 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_995 <= 32'h0;
    end else begin
      if (11'h3e3 == _T_12323) begin
        mem_995 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_996 <= 32'h0;
    end else begin
      if (11'h3e4 == _T_12323) begin
        mem_996 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_997 <= 32'h0;
    end else begin
      if (11'h3e5 == _T_12323) begin
        mem_997 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_998 <= 32'h0;
    end else begin
      if (11'h3e6 == _T_12323) begin
        mem_998 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_999 <= 32'h0;
    end else begin
      if (11'h3e7 == _T_12323) begin
        mem_999 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1000 <= 32'h0;
    end else begin
      if (11'h3e8 == _T_12323) begin
        mem_1000 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1001 <= 32'h0;
    end else begin
      if (11'h3e9 == _T_12323) begin
        mem_1001 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1002 <= 32'h0;
    end else begin
      if (11'h3ea == _T_12323) begin
        mem_1002 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1003 <= 32'h0;
    end else begin
      if (11'h3eb == _T_12323) begin
        mem_1003 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1004 <= 32'h0;
    end else begin
      if (11'h3ec == _T_12323) begin
        mem_1004 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1005 <= 32'h0;
    end else begin
      if (11'h3ed == _T_12323) begin
        mem_1005 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1006 <= 32'h0;
    end else begin
      if (11'h3ee == _T_12323) begin
        mem_1006 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1007 <= 32'h0;
    end else begin
      if (11'h3ef == _T_12323) begin
        mem_1007 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1008 <= 32'h0;
    end else begin
      if (11'h3f0 == _T_12323) begin
        mem_1008 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1009 <= 32'h0;
    end else begin
      if (11'h3f1 == _T_12323) begin
        mem_1009 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1010 <= 32'h0;
    end else begin
      if (11'h3f2 == _T_12323) begin
        mem_1010 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1011 <= 32'h0;
    end else begin
      if (11'h3f3 == _T_12323) begin
        mem_1011 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1012 <= 32'h0;
    end else begin
      if (11'h3f4 == _T_12323) begin
        mem_1012 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1013 <= 32'h0;
    end else begin
      if (11'h3f5 == _T_12323) begin
        mem_1013 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1014 <= 32'h0;
    end else begin
      if (11'h3f6 == _T_12323) begin
        mem_1014 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1015 <= 32'h0;
    end else begin
      if (11'h3f7 == _T_12323) begin
        mem_1015 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1016 <= 32'h0;
    end else begin
      if (11'h3f8 == _T_12323) begin
        mem_1016 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1017 <= 32'h0;
    end else begin
      if (11'h3f9 == _T_12323) begin
        mem_1017 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1018 <= 32'h0;
    end else begin
      if (11'h3fa == _T_12323) begin
        mem_1018 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1019 <= 32'h0;
    end else begin
      if (11'h3fb == _T_12323) begin
        mem_1019 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1020 <= 32'h0;
    end else begin
      if (11'h3fc == _T_12323) begin
        mem_1020 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1021 <= 32'h0;
    end else begin
      if (11'h3fd == _T_12323) begin
        mem_1021 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1022 <= 32'h0;
    end else begin
      if (11'h3fe == _T_12323) begin
        mem_1022 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1023 <= 32'h0;
    end else begin
      if (11'h3ff == _T_12323) begin
        mem_1023 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1024 <= 32'h0;
    end else begin
      if (11'h400 == _T_12323) begin
        mem_1024 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1025 <= 32'h0;
    end else begin
      if (11'h401 == _T_12323) begin
        mem_1025 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1026 <= 32'h0;
    end else begin
      if (11'h402 == _T_12323) begin
        mem_1026 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1027 <= 32'h0;
    end else begin
      if (11'h403 == _T_12323) begin
        mem_1027 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1028 <= 32'h0;
    end else begin
      if (11'h404 == _T_12323) begin
        mem_1028 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1029 <= 32'h0;
    end else begin
      if (11'h405 == _T_12323) begin
        mem_1029 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1030 <= 32'h0;
    end else begin
      if (11'h406 == _T_12323) begin
        mem_1030 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1031 <= 32'h0;
    end else begin
      if (11'h407 == _T_12323) begin
        mem_1031 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1032 <= 32'h0;
    end else begin
      if (11'h408 == _T_12323) begin
        mem_1032 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1033 <= 32'h0;
    end else begin
      if (11'h409 == _T_12323) begin
        mem_1033 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1034 <= 32'h0;
    end else begin
      if (11'h40a == _T_12323) begin
        mem_1034 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1035 <= 32'h0;
    end else begin
      if (11'h40b == _T_12323) begin
        mem_1035 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1036 <= 32'h0;
    end else begin
      if (11'h40c == _T_12323) begin
        mem_1036 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1037 <= 32'h0;
    end else begin
      if (11'h40d == _T_12323) begin
        mem_1037 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1038 <= 32'h0;
    end else begin
      if (11'h40e == _T_12323) begin
        mem_1038 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1039 <= 32'h0;
    end else begin
      if (11'h40f == _T_12323) begin
        mem_1039 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1040 <= 32'h0;
    end else begin
      if (11'h410 == _T_12323) begin
        mem_1040 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1041 <= 32'h0;
    end else begin
      if (11'h411 == _T_12323) begin
        mem_1041 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1042 <= 32'h0;
    end else begin
      if (11'h412 == _T_12323) begin
        mem_1042 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1043 <= 32'h0;
    end else begin
      if (11'h413 == _T_12323) begin
        mem_1043 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1044 <= 32'h0;
    end else begin
      if (11'h414 == _T_12323) begin
        mem_1044 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1045 <= 32'h0;
    end else begin
      if (11'h415 == _T_12323) begin
        mem_1045 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1046 <= 32'h0;
    end else begin
      if (11'h416 == _T_12323) begin
        mem_1046 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1047 <= 32'h0;
    end else begin
      if (11'h417 == _T_12323) begin
        mem_1047 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1048 <= 32'h0;
    end else begin
      if (11'h418 == _T_12323) begin
        mem_1048 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1049 <= 32'h0;
    end else begin
      if (11'h419 == _T_12323) begin
        mem_1049 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1050 <= 32'h0;
    end else begin
      if (11'h41a == _T_12323) begin
        mem_1050 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1051 <= 32'h0;
    end else begin
      if (11'h41b == _T_12323) begin
        mem_1051 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1052 <= 32'h0;
    end else begin
      if (11'h41c == _T_12323) begin
        mem_1052 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1053 <= 32'h0;
    end else begin
      if (11'h41d == _T_12323) begin
        mem_1053 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1054 <= 32'h0;
    end else begin
      if (11'h41e == _T_12323) begin
        mem_1054 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1055 <= 32'h0;
    end else begin
      if (11'h41f == _T_12323) begin
        mem_1055 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1056 <= 32'h0;
    end else begin
      if (11'h420 == _T_12323) begin
        mem_1056 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1057 <= 32'h0;
    end else begin
      if (11'h421 == _T_12323) begin
        mem_1057 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1058 <= 32'h0;
    end else begin
      if (11'h422 == _T_12323) begin
        mem_1058 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1059 <= 32'h0;
    end else begin
      if (11'h423 == _T_12323) begin
        mem_1059 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1060 <= 32'h0;
    end else begin
      if (11'h424 == _T_12323) begin
        mem_1060 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1061 <= 32'h0;
    end else begin
      if (11'h425 == _T_12323) begin
        mem_1061 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1062 <= 32'h0;
    end else begin
      if (11'h426 == _T_12323) begin
        mem_1062 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1063 <= 32'h0;
    end else begin
      if (11'h427 == _T_12323) begin
        mem_1063 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1064 <= 32'h0;
    end else begin
      if (11'h428 == _T_12323) begin
        mem_1064 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1065 <= 32'h0;
    end else begin
      if (11'h429 == _T_12323) begin
        mem_1065 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1066 <= 32'h0;
    end else begin
      if (11'h42a == _T_12323) begin
        mem_1066 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1067 <= 32'h0;
    end else begin
      if (11'h42b == _T_12323) begin
        mem_1067 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1068 <= 32'h0;
    end else begin
      if (11'h42c == _T_12323) begin
        mem_1068 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1069 <= 32'h0;
    end else begin
      if (11'h42d == _T_12323) begin
        mem_1069 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1070 <= 32'h0;
    end else begin
      if (11'h42e == _T_12323) begin
        mem_1070 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1071 <= 32'h0;
    end else begin
      if (11'h42f == _T_12323) begin
        mem_1071 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1072 <= 32'h0;
    end else begin
      if (11'h430 == _T_12323) begin
        mem_1072 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1073 <= 32'h0;
    end else begin
      if (11'h431 == _T_12323) begin
        mem_1073 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1074 <= 32'h0;
    end else begin
      if (11'h432 == _T_12323) begin
        mem_1074 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1075 <= 32'h0;
    end else begin
      if (11'h433 == _T_12323) begin
        mem_1075 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1076 <= 32'h0;
    end else begin
      if (11'h434 == _T_12323) begin
        mem_1076 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1077 <= 32'h0;
    end else begin
      if (11'h435 == _T_12323) begin
        mem_1077 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1078 <= 32'h0;
    end else begin
      if (11'h436 == _T_12323) begin
        mem_1078 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1079 <= 32'h0;
    end else begin
      if (11'h437 == _T_12323) begin
        mem_1079 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1080 <= 32'h0;
    end else begin
      if (11'h438 == _T_12323) begin
        mem_1080 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1081 <= 32'h0;
    end else begin
      if (11'h439 == _T_12323) begin
        mem_1081 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1082 <= 32'h0;
    end else begin
      if (11'h43a == _T_12323) begin
        mem_1082 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1083 <= 32'h0;
    end else begin
      if (11'h43b == _T_12323) begin
        mem_1083 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1084 <= 32'h0;
    end else begin
      if (11'h43c == _T_12323) begin
        mem_1084 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1085 <= 32'h0;
    end else begin
      if (11'h43d == _T_12323) begin
        mem_1085 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1086 <= 32'h0;
    end else begin
      if (11'h43e == _T_12323) begin
        mem_1086 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1087 <= 32'h0;
    end else begin
      if (11'h43f == _T_12323) begin
        mem_1087 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1088 <= 32'h0;
    end else begin
      if (11'h440 == _T_12323) begin
        mem_1088 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1089 <= 32'h0;
    end else begin
      if (11'h441 == _T_12323) begin
        mem_1089 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1090 <= 32'h0;
    end else begin
      if (11'h442 == _T_12323) begin
        mem_1090 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1091 <= 32'h0;
    end else begin
      if (11'h443 == _T_12323) begin
        mem_1091 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1092 <= 32'h0;
    end else begin
      if (11'h444 == _T_12323) begin
        mem_1092 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1093 <= 32'h0;
    end else begin
      if (11'h445 == _T_12323) begin
        mem_1093 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1094 <= 32'h0;
    end else begin
      if (11'h446 == _T_12323) begin
        mem_1094 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1095 <= 32'h0;
    end else begin
      if (11'h447 == _T_12323) begin
        mem_1095 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1096 <= 32'h0;
    end else begin
      if (11'h448 == _T_12323) begin
        mem_1096 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1097 <= 32'h0;
    end else begin
      if (11'h449 == _T_12323) begin
        mem_1097 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1098 <= 32'h0;
    end else begin
      if (11'h44a == _T_12323) begin
        mem_1098 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1099 <= 32'h0;
    end else begin
      if (11'h44b == _T_12323) begin
        mem_1099 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1100 <= 32'h0;
    end else begin
      if (11'h44c == _T_12323) begin
        mem_1100 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1101 <= 32'h0;
    end else begin
      if (11'h44d == _T_12323) begin
        mem_1101 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1102 <= 32'h0;
    end else begin
      if (11'h44e == _T_12323) begin
        mem_1102 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1103 <= 32'h0;
    end else begin
      if (11'h44f == _T_12323) begin
        mem_1103 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1104 <= 32'h0;
    end else begin
      if (11'h450 == _T_12323) begin
        mem_1104 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1105 <= 32'h0;
    end else begin
      if (11'h451 == _T_12323) begin
        mem_1105 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1106 <= 32'h0;
    end else begin
      if (11'h452 == _T_12323) begin
        mem_1106 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1107 <= 32'h0;
    end else begin
      if (11'h453 == _T_12323) begin
        mem_1107 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1108 <= 32'h0;
    end else begin
      if (11'h454 == _T_12323) begin
        mem_1108 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1109 <= 32'h0;
    end else begin
      if (11'h455 == _T_12323) begin
        mem_1109 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1110 <= 32'h0;
    end else begin
      if (11'h456 == _T_12323) begin
        mem_1110 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1111 <= 32'h0;
    end else begin
      if (11'h457 == _T_12323) begin
        mem_1111 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1112 <= 32'h0;
    end else begin
      if (11'h458 == _T_12323) begin
        mem_1112 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1113 <= 32'h0;
    end else begin
      if (11'h459 == _T_12323) begin
        mem_1113 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1114 <= 32'h0;
    end else begin
      if (11'h45a == _T_12323) begin
        mem_1114 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1115 <= 32'h0;
    end else begin
      if (11'h45b == _T_12323) begin
        mem_1115 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1116 <= 32'h0;
    end else begin
      if (11'h45c == _T_12323) begin
        mem_1116 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1117 <= 32'h0;
    end else begin
      if (11'h45d == _T_12323) begin
        mem_1117 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1118 <= 32'h0;
    end else begin
      if (11'h45e == _T_12323) begin
        mem_1118 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1119 <= 32'h0;
    end else begin
      if (11'h45f == _T_12323) begin
        mem_1119 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1120 <= 32'h0;
    end else begin
      if (11'h460 == _T_12323) begin
        mem_1120 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1121 <= 32'h0;
    end else begin
      if (11'h461 == _T_12323) begin
        mem_1121 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1122 <= 32'h0;
    end else begin
      if (11'h462 == _T_12323) begin
        mem_1122 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1123 <= 32'h0;
    end else begin
      if (11'h463 == _T_12323) begin
        mem_1123 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1124 <= 32'h0;
    end else begin
      if (11'h464 == _T_12323) begin
        mem_1124 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1125 <= 32'h0;
    end else begin
      if (11'h465 == _T_12323) begin
        mem_1125 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1126 <= 32'h0;
    end else begin
      if (11'h466 == _T_12323) begin
        mem_1126 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1127 <= 32'h0;
    end else begin
      if (11'h467 == _T_12323) begin
        mem_1127 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1128 <= 32'h0;
    end else begin
      if (11'h468 == _T_12323) begin
        mem_1128 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1129 <= 32'h0;
    end else begin
      if (11'h469 == _T_12323) begin
        mem_1129 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1130 <= 32'h0;
    end else begin
      if (11'h46a == _T_12323) begin
        mem_1130 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1131 <= 32'h0;
    end else begin
      if (11'h46b == _T_12323) begin
        mem_1131 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1132 <= 32'h0;
    end else begin
      if (11'h46c == _T_12323) begin
        mem_1132 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1133 <= 32'h0;
    end else begin
      if (11'h46d == _T_12323) begin
        mem_1133 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1134 <= 32'h0;
    end else begin
      if (11'h46e == _T_12323) begin
        mem_1134 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1135 <= 32'h0;
    end else begin
      if (11'h46f == _T_12323) begin
        mem_1135 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1136 <= 32'h0;
    end else begin
      if (11'h470 == _T_12323) begin
        mem_1136 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1137 <= 32'h0;
    end else begin
      if (11'h471 == _T_12323) begin
        mem_1137 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1138 <= 32'h0;
    end else begin
      if (11'h472 == _T_12323) begin
        mem_1138 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1139 <= 32'h0;
    end else begin
      if (11'h473 == _T_12323) begin
        mem_1139 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1140 <= 32'h0;
    end else begin
      if (11'h474 == _T_12323) begin
        mem_1140 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1141 <= 32'h0;
    end else begin
      if (11'h475 == _T_12323) begin
        mem_1141 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1142 <= 32'h0;
    end else begin
      if (11'h476 == _T_12323) begin
        mem_1142 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1143 <= 32'h0;
    end else begin
      if (11'h477 == _T_12323) begin
        mem_1143 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1144 <= 32'h0;
    end else begin
      if (11'h478 == _T_12323) begin
        mem_1144 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1145 <= 32'h0;
    end else begin
      if (11'h479 == _T_12323) begin
        mem_1145 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1146 <= 32'h0;
    end else begin
      if (11'h47a == _T_12323) begin
        mem_1146 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1147 <= 32'h0;
    end else begin
      if (11'h47b == _T_12323) begin
        mem_1147 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1148 <= 32'h0;
    end else begin
      if (11'h47c == _T_12323) begin
        mem_1148 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1149 <= 32'h0;
    end else begin
      if (11'h47d == _T_12323) begin
        mem_1149 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1150 <= 32'h0;
    end else begin
      if (11'h47e == _T_12323) begin
        mem_1150 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1151 <= 32'h0;
    end else begin
      if (11'h47f == _T_12323) begin
        mem_1151 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1152 <= 32'h0;
    end else begin
      if (11'h480 == _T_12323) begin
        mem_1152 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1153 <= 32'h0;
    end else begin
      if (11'h481 == _T_12323) begin
        mem_1153 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1154 <= 32'h0;
    end else begin
      if (11'h482 == _T_12323) begin
        mem_1154 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1155 <= 32'h0;
    end else begin
      if (11'h483 == _T_12323) begin
        mem_1155 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1156 <= 32'h0;
    end else begin
      if (11'h484 == _T_12323) begin
        mem_1156 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1157 <= 32'h0;
    end else begin
      if (11'h485 == _T_12323) begin
        mem_1157 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1158 <= 32'h0;
    end else begin
      if (11'h486 == _T_12323) begin
        mem_1158 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1159 <= 32'h0;
    end else begin
      if (11'h487 == _T_12323) begin
        mem_1159 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1160 <= 32'h0;
    end else begin
      if (11'h488 == _T_12323) begin
        mem_1160 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1161 <= 32'h0;
    end else begin
      if (11'h489 == _T_12323) begin
        mem_1161 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1162 <= 32'h0;
    end else begin
      if (11'h48a == _T_12323) begin
        mem_1162 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1163 <= 32'h0;
    end else begin
      if (11'h48b == _T_12323) begin
        mem_1163 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1164 <= 32'h0;
    end else begin
      if (11'h48c == _T_12323) begin
        mem_1164 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1165 <= 32'h0;
    end else begin
      if (11'h48d == _T_12323) begin
        mem_1165 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1166 <= 32'h0;
    end else begin
      if (11'h48e == _T_12323) begin
        mem_1166 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1167 <= 32'h0;
    end else begin
      if (11'h48f == _T_12323) begin
        mem_1167 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1168 <= 32'h0;
    end else begin
      if (11'h490 == _T_12323) begin
        mem_1168 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1169 <= 32'h0;
    end else begin
      if (11'h491 == _T_12323) begin
        mem_1169 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1170 <= 32'h0;
    end else begin
      if (11'h492 == _T_12323) begin
        mem_1170 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1171 <= 32'h0;
    end else begin
      if (11'h493 == _T_12323) begin
        mem_1171 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1172 <= 32'h0;
    end else begin
      if (11'h494 == _T_12323) begin
        mem_1172 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1173 <= 32'h0;
    end else begin
      if (11'h495 == _T_12323) begin
        mem_1173 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1174 <= 32'h0;
    end else begin
      if (11'h496 == _T_12323) begin
        mem_1174 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1175 <= 32'h0;
    end else begin
      if (11'h497 == _T_12323) begin
        mem_1175 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1176 <= 32'h0;
    end else begin
      if (11'h498 == _T_12323) begin
        mem_1176 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1177 <= 32'h0;
    end else begin
      if (11'h499 == _T_12323) begin
        mem_1177 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1178 <= 32'h0;
    end else begin
      if (11'h49a == _T_12323) begin
        mem_1178 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1179 <= 32'h0;
    end else begin
      if (11'h49b == _T_12323) begin
        mem_1179 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1180 <= 32'h0;
    end else begin
      if (11'h49c == _T_12323) begin
        mem_1180 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1181 <= 32'h0;
    end else begin
      if (11'h49d == _T_12323) begin
        mem_1181 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1182 <= 32'h0;
    end else begin
      if (11'h49e == _T_12323) begin
        mem_1182 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1183 <= 32'h0;
    end else begin
      if (11'h49f == _T_12323) begin
        mem_1183 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1184 <= 32'h0;
    end else begin
      if (11'h4a0 == _T_12323) begin
        mem_1184 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1185 <= 32'h0;
    end else begin
      if (11'h4a1 == _T_12323) begin
        mem_1185 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1186 <= 32'h0;
    end else begin
      if (11'h4a2 == _T_12323) begin
        mem_1186 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1187 <= 32'h0;
    end else begin
      if (11'h4a3 == _T_12323) begin
        mem_1187 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1188 <= 32'h0;
    end else begin
      if (11'h4a4 == _T_12323) begin
        mem_1188 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1189 <= 32'h0;
    end else begin
      if (11'h4a5 == _T_12323) begin
        mem_1189 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1190 <= 32'h0;
    end else begin
      if (11'h4a6 == _T_12323) begin
        mem_1190 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1191 <= 32'h0;
    end else begin
      if (11'h4a7 == _T_12323) begin
        mem_1191 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1192 <= 32'h0;
    end else begin
      if (11'h4a8 == _T_12323) begin
        mem_1192 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1193 <= 32'h0;
    end else begin
      if (11'h4a9 == _T_12323) begin
        mem_1193 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1194 <= 32'h0;
    end else begin
      if (11'h4aa == _T_12323) begin
        mem_1194 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1195 <= 32'h0;
    end else begin
      if (11'h4ab == _T_12323) begin
        mem_1195 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1196 <= 32'h0;
    end else begin
      if (11'h4ac == _T_12323) begin
        mem_1196 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1197 <= 32'h0;
    end else begin
      if (11'h4ad == _T_12323) begin
        mem_1197 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1198 <= 32'h0;
    end else begin
      if (11'h4ae == _T_12323) begin
        mem_1198 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1199 <= 32'h0;
    end else begin
      if (11'h4af == _T_12323) begin
        mem_1199 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1200 <= 32'h0;
    end else begin
      if (11'h4b0 == _T_12323) begin
        mem_1200 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1201 <= 32'h0;
    end else begin
      if (11'h4b1 == _T_12323) begin
        mem_1201 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1202 <= 32'h0;
    end else begin
      if (11'h4b2 == _T_12323) begin
        mem_1202 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1203 <= 32'h0;
    end else begin
      if (11'h4b3 == _T_12323) begin
        mem_1203 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1204 <= 32'h0;
    end else begin
      if (11'h4b4 == _T_12323) begin
        mem_1204 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1205 <= 32'h0;
    end else begin
      if (11'h4b5 == _T_12323) begin
        mem_1205 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1206 <= 32'h0;
    end else begin
      if (11'h4b6 == _T_12323) begin
        mem_1206 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1207 <= 32'h0;
    end else begin
      if (11'h4b7 == _T_12323) begin
        mem_1207 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1208 <= 32'h0;
    end else begin
      if (11'h4b8 == _T_12323) begin
        mem_1208 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1209 <= 32'h0;
    end else begin
      if (11'h4b9 == _T_12323) begin
        mem_1209 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1210 <= 32'h0;
    end else begin
      if (11'h4ba == _T_12323) begin
        mem_1210 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1211 <= 32'h0;
    end else begin
      if (11'h4bb == _T_12323) begin
        mem_1211 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1212 <= 32'h0;
    end else begin
      if (11'h4bc == _T_12323) begin
        mem_1212 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1213 <= 32'h0;
    end else begin
      if (11'h4bd == _T_12323) begin
        mem_1213 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1214 <= 32'h0;
    end else begin
      if (11'h4be == _T_12323) begin
        mem_1214 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1215 <= 32'h0;
    end else begin
      if (11'h4bf == _T_12323) begin
        mem_1215 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1216 <= 32'h0;
    end else begin
      if (11'h4c0 == _T_12323) begin
        mem_1216 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1217 <= 32'h0;
    end else begin
      if (11'h4c1 == _T_12323) begin
        mem_1217 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1218 <= 32'h0;
    end else begin
      if (11'h4c2 == _T_12323) begin
        mem_1218 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1219 <= 32'h0;
    end else begin
      if (11'h4c3 == _T_12323) begin
        mem_1219 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1220 <= 32'h0;
    end else begin
      if (11'h4c4 == _T_12323) begin
        mem_1220 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1221 <= 32'h0;
    end else begin
      if (11'h4c5 == _T_12323) begin
        mem_1221 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1222 <= 32'h0;
    end else begin
      if (11'h4c6 == _T_12323) begin
        mem_1222 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1223 <= 32'h0;
    end else begin
      if (11'h4c7 == _T_12323) begin
        mem_1223 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1224 <= 32'h0;
    end else begin
      if (11'h4c8 == _T_12323) begin
        mem_1224 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1225 <= 32'h0;
    end else begin
      if (11'h4c9 == _T_12323) begin
        mem_1225 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1226 <= 32'h0;
    end else begin
      if (11'h4ca == _T_12323) begin
        mem_1226 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1227 <= 32'h0;
    end else begin
      if (11'h4cb == _T_12323) begin
        mem_1227 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1228 <= 32'h0;
    end else begin
      if (11'h4cc == _T_12323) begin
        mem_1228 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1229 <= 32'h0;
    end else begin
      if (11'h4cd == _T_12323) begin
        mem_1229 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1230 <= 32'h0;
    end else begin
      if (11'h4ce == _T_12323) begin
        mem_1230 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1231 <= 32'h0;
    end else begin
      if (11'h4cf == _T_12323) begin
        mem_1231 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1232 <= 32'h0;
    end else begin
      if (11'h4d0 == _T_12323) begin
        mem_1232 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1233 <= 32'h0;
    end else begin
      if (11'h4d1 == _T_12323) begin
        mem_1233 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1234 <= 32'h0;
    end else begin
      if (11'h4d2 == _T_12323) begin
        mem_1234 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1235 <= 32'h0;
    end else begin
      if (11'h4d3 == _T_12323) begin
        mem_1235 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1236 <= 32'h0;
    end else begin
      if (11'h4d4 == _T_12323) begin
        mem_1236 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1237 <= 32'h0;
    end else begin
      if (11'h4d5 == _T_12323) begin
        mem_1237 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1238 <= 32'h0;
    end else begin
      if (11'h4d6 == _T_12323) begin
        mem_1238 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1239 <= 32'h0;
    end else begin
      if (11'h4d7 == _T_12323) begin
        mem_1239 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1240 <= 32'h0;
    end else begin
      if (11'h4d8 == _T_12323) begin
        mem_1240 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1241 <= 32'h0;
    end else begin
      if (11'h4d9 == _T_12323) begin
        mem_1241 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1242 <= 32'h0;
    end else begin
      if (11'h4da == _T_12323) begin
        mem_1242 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1243 <= 32'h0;
    end else begin
      if (11'h4db == _T_12323) begin
        mem_1243 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1244 <= 32'h0;
    end else begin
      if (11'h4dc == _T_12323) begin
        mem_1244 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1245 <= 32'h0;
    end else begin
      if (11'h4dd == _T_12323) begin
        mem_1245 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1246 <= 32'h0;
    end else begin
      if (11'h4de == _T_12323) begin
        mem_1246 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1247 <= 32'h0;
    end else begin
      if (11'h4df == _T_12323) begin
        mem_1247 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1248 <= 32'h0;
    end else begin
      if (11'h4e0 == _T_12323) begin
        mem_1248 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1249 <= 32'h0;
    end else begin
      if (11'h4e1 == _T_12323) begin
        mem_1249 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1250 <= 32'h0;
    end else begin
      if (11'h4e2 == _T_12323) begin
        mem_1250 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1251 <= 32'h0;
    end else begin
      if (11'h4e3 == _T_12323) begin
        mem_1251 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1252 <= 32'h0;
    end else begin
      if (11'h4e4 == _T_12323) begin
        mem_1252 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1253 <= 32'h0;
    end else begin
      if (11'h4e5 == _T_12323) begin
        mem_1253 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1254 <= 32'h0;
    end else begin
      if (11'h4e6 == _T_12323) begin
        mem_1254 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1255 <= 32'h0;
    end else begin
      if (11'h4e7 == _T_12323) begin
        mem_1255 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1256 <= 32'h0;
    end else begin
      if (11'h4e8 == _T_12323) begin
        mem_1256 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1257 <= 32'h0;
    end else begin
      if (11'h4e9 == _T_12323) begin
        mem_1257 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1258 <= 32'h0;
    end else begin
      if (11'h4ea == _T_12323) begin
        mem_1258 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1259 <= 32'h0;
    end else begin
      if (11'h4eb == _T_12323) begin
        mem_1259 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1260 <= 32'h0;
    end else begin
      if (11'h4ec == _T_12323) begin
        mem_1260 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1261 <= 32'h0;
    end else begin
      if (11'h4ed == _T_12323) begin
        mem_1261 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1262 <= 32'h0;
    end else begin
      if (11'h4ee == _T_12323) begin
        mem_1262 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1263 <= 32'h0;
    end else begin
      if (11'h4ef == _T_12323) begin
        mem_1263 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1264 <= 32'h0;
    end else begin
      if (11'h4f0 == _T_12323) begin
        mem_1264 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1265 <= 32'h0;
    end else begin
      if (11'h4f1 == _T_12323) begin
        mem_1265 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1266 <= 32'h0;
    end else begin
      if (11'h4f2 == _T_12323) begin
        mem_1266 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1267 <= 32'h0;
    end else begin
      if (11'h4f3 == _T_12323) begin
        mem_1267 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1268 <= 32'h0;
    end else begin
      if (11'h4f4 == _T_12323) begin
        mem_1268 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1269 <= 32'h0;
    end else begin
      if (11'h4f5 == _T_12323) begin
        mem_1269 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1270 <= 32'h0;
    end else begin
      if (11'h4f6 == _T_12323) begin
        mem_1270 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1271 <= 32'h0;
    end else begin
      if (11'h4f7 == _T_12323) begin
        mem_1271 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1272 <= 32'h0;
    end else begin
      if (11'h4f8 == _T_12323) begin
        mem_1272 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1273 <= 32'h0;
    end else begin
      if (11'h4f9 == _T_12323) begin
        mem_1273 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1274 <= 32'h0;
    end else begin
      if (11'h4fa == _T_12323) begin
        mem_1274 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1275 <= 32'h0;
    end else begin
      if (11'h4fb == _T_12323) begin
        mem_1275 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1276 <= 32'h0;
    end else begin
      if (11'h4fc == _T_12323) begin
        mem_1276 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1277 <= 32'h0;
    end else begin
      if (11'h4fd == _T_12323) begin
        mem_1277 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1278 <= 32'h0;
    end else begin
      if (11'h4fe == _T_12323) begin
        mem_1278 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1279 <= 32'h0;
    end else begin
      if (11'h4ff == _T_12323) begin
        mem_1279 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1280 <= 32'h0;
    end else begin
      if (11'h500 == _T_12323) begin
        mem_1280 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1281 <= 32'h0;
    end else begin
      if (11'h501 == _T_12323) begin
        mem_1281 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1282 <= 32'h0;
    end else begin
      if (11'h502 == _T_12323) begin
        mem_1282 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1283 <= 32'h0;
    end else begin
      if (11'h503 == _T_12323) begin
        mem_1283 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1284 <= 32'h0;
    end else begin
      if (11'h504 == _T_12323) begin
        mem_1284 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1285 <= 32'h0;
    end else begin
      if (11'h505 == _T_12323) begin
        mem_1285 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1286 <= 32'h0;
    end else begin
      if (11'h506 == _T_12323) begin
        mem_1286 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1287 <= 32'h0;
    end else begin
      if (11'h507 == _T_12323) begin
        mem_1287 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1288 <= 32'h0;
    end else begin
      if (11'h508 == _T_12323) begin
        mem_1288 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1289 <= 32'h0;
    end else begin
      if (11'h509 == _T_12323) begin
        mem_1289 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1290 <= 32'h0;
    end else begin
      if (11'h50a == _T_12323) begin
        mem_1290 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1291 <= 32'h0;
    end else begin
      if (11'h50b == _T_12323) begin
        mem_1291 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1292 <= 32'h0;
    end else begin
      if (11'h50c == _T_12323) begin
        mem_1292 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1293 <= 32'h0;
    end else begin
      if (11'h50d == _T_12323) begin
        mem_1293 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1294 <= 32'h0;
    end else begin
      if (11'h50e == _T_12323) begin
        mem_1294 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1295 <= 32'h0;
    end else begin
      if (11'h50f == _T_12323) begin
        mem_1295 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1296 <= 32'h0;
    end else begin
      if (11'h510 == _T_12323) begin
        mem_1296 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1297 <= 32'h0;
    end else begin
      if (11'h511 == _T_12323) begin
        mem_1297 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1298 <= 32'h0;
    end else begin
      if (11'h512 == _T_12323) begin
        mem_1298 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1299 <= 32'h0;
    end else begin
      if (11'h513 == _T_12323) begin
        mem_1299 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1300 <= 32'h0;
    end else begin
      if (11'h514 == _T_12323) begin
        mem_1300 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1301 <= 32'h0;
    end else begin
      if (11'h515 == _T_12323) begin
        mem_1301 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1302 <= 32'h0;
    end else begin
      if (11'h516 == _T_12323) begin
        mem_1302 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1303 <= 32'h0;
    end else begin
      if (11'h517 == _T_12323) begin
        mem_1303 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1304 <= 32'h0;
    end else begin
      if (11'h518 == _T_12323) begin
        mem_1304 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1305 <= 32'h0;
    end else begin
      if (11'h519 == _T_12323) begin
        mem_1305 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1306 <= 32'h0;
    end else begin
      if (11'h51a == _T_12323) begin
        mem_1306 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1307 <= 32'h0;
    end else begin
      if (11'h51b == _T_12323) begin
        mem_1307 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1308 <= 32'h0;
    end else begin
      if (11'h51c == _T_12323) begin
        mem_1308 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1309 <= 32'h0;
    end else begin
      if (11'h51d == _T_12323) begin
        mem_1309 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1310 <= 32'h0;
    end else begin
      if (11'h51e == _T_12323) begin
        mem_1310 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1311 <= 32'h0;
    end else begin
      if (11'h51f == _T_12323) begin
        mem_1311 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1312 <= 32'h0;
    end else begin
      if (11'h520 == _T_12323) begin
        mem_1312 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1313 <= 32'h0;
    end else begin
      if (11'h521 == _T_12323) begin
        mem_1313 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1314 <= 32'h0;
    end else begin
      if (11'h522 == _T_12323) begin
        mem_1314 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1315 <= 32'h0;
    end else begin
      if (11'h523 == _T_12323) begin
        mem_1315 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1316 <= 32'h0;
    end else begin
      if (11'h524 == _T_12323) begin
        mem_1316 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1317 <= 32'h0;
    end else begin
      if (11'h525 == _T_12323) begin
        mem_1317 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1318 <= 32'h0;
    end else begin
      if (11'h526 == _T_12323) begin
        mem_1318 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1319 <= 32'h0;
    end else begin
      if (11'h527 == _T_12323) begin
        mem_1319 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1320 <= 32'h0;
    end else begin
      if (11'h528 == _T_12323) begin
        mem_1320 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1321 <= 32'h0;
    end else begin
      if (11'h529 == _T_12323) begin
        mem_1321 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1322 <= 32'h0;
    end else begin
      if (11'h52a == _T_12323) begin
        mem_1322 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1323 <= 32'h0;
    end else begin
      if (11'h52b == _T_12323) begin
        mem_1323 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1324 <= 32'h0;
    end else begin
      if (11'h52c == _T_12323) begin
        mem_1324 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1325 <= 32'h0;
    end else begin
      if (11'h52d == _T_12323) begin
        mem_1325 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1326 <= 32'h0;
    end else begin
      if (11'h52e == _T_12323) begin
        mem_1326 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1327 <= 32'h0;
    end else begin
      if (11'h52f == _T_12323) begin
        mem_1327 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1328 <= 32'h0;
    end else begin
      if (11'h530 == _T_12323) begin
        mem_1328 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1329 <= 32'h0;
    end else begin
      if (11'h531 == _T_12323) begin
        mem_1329 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1330 <= 32'h0;
    end else begin
      if (11'h532 == _T_12323) begin
        mem_1330 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1331 <= 32'h0;
    end else begin
      if (11'h533 == _T_12323) begin
        mem_1331 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1332 <= 32'h0;
    end else begin
      if (11'h534 == _T_12323) begin
        mem_1332 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1333 <= 32'h0;
    end else begin
      if (11'h535 == _T_12323) begin
        mem_1333 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1334 <= 32'h0;
    end else begin
      if (11'h536 == _T_12323) begin
        mem_1334 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1335 <= 32'h0;
    end else begin
      if (11'h537 == _T_12323) begin
        mem_1335 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1336 <= 32'h0;
    end else begin
      if (11'h538 == _T_12323) begin
        mem_1336 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1337 <= 32'h0;
    end else begin
      if (11'h539 == _T_12323) begin
        mem_1337 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1338 <= 32'h0;
    end else begin
      if (11'h53a == _T_12323) begin
        mem_1338 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1339 <= 32'h0;
    end else begin
      if (11'h53b == _T_12323) begin
        mem_1339 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1340 <= 32'h0;
    end else begin
      if (11'h53c == _T_12323) begin
        mem_1340 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1341 <= 32'h0;
    end else begin
      if (11'h53d == _T_12323) begin
        mem_1341 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1342 <= 32'h0;
    end else begin
      if (11'h53e == _T_12323) begin
        mem_1342 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1343 <= 32'h0;
    end else begin
      if (11'h53f == _T_12323) begin
        mem_1343 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1344 <= 32'h0;
    end else begin
      if (11'h540 == _T_12323) begin
        mem_1344 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1345 <= 32'h0;
    end else begin
      if (11'h541 == _T_12323) begin
        mem_1345 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1346 <= 32'h0;
    end else begin
      if (11'h542 == _T_12323) begin
        mem_1346 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1347 <= 32'h0;
    end else begin
      if (11'h543 == _T_12323) begin
        mem_1347 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1348 <= 32'h0;
    end else begin
      if (11'h544 == _T_12323) begin
        mem_1348 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1349 <= 32'h0;
    end else begin
      if (11'h545 == _T_12323) begin
        mem_1349 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1350 <= 32'h0;
    end else begin
      if (11'h546 == _T_12323) begin
        mem_1350 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1351 <= 32'h0;
    end else begin
      if (11'h547 == _T_12323) begin
        mem_1351 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1352 <= 32'h0;
    end else begin
      if (11'h548 == _T_12323) begin
        mem_1352 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1353 <= 32'h0;
    end else begin
      if (11'h549 == _T_12323) begin
        mem_1353 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1354 <= 32'h0;
    end else begin
      if (11'h54a == _T_12323) begin
        mem_1354 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1355 <= 32'h0;
    end else begin
      if (11'h54b == _T_12323) begin
        mem_1355 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1356 <= 32'h0;
    end else begin
      if (11'h54c == _T_12323) begin
        mem_1356 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1357 <= 32'h0;
    end else begin
      if (11'h54d == _T_12323) begin
        mem_1357 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1358 <= 32'h0;
    end else begin
      if (11'h54e == _T_12323) begin
        mem_1358 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1359 <= 32'h0;
    end else begin
      if (11'h54f == _T_12323) begin
        mem_1359 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1360 <= 32'h0;
    end else begin
      if (11'h550 == _T_12323) begin
        mem_1360 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1361 <= 32'h0;
    end else begin
      if (11'h551 == _T_12323) begin
        mem_1361 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1362 <= 32'h0;
    end else begin
      if (11'h552 == _T_12323) begin
        mem_1362 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1363 <= 32'h0;
    end else begin
      if (11'h553 == _T_12323) begin
        mem_1363 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1364 <= 32'h0;
    end else begin
      if (11'h554 == _T_12323) begin
        mem_1364 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1365 <= 32'h0;
    end else begin
      if (11'h555 == _T_12323) begin
        mem_1365 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1366 <= 32'h0;
    end else begin
      if (11'h556 == _T_12323) begin
        mem_1366 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1367 <= 32'h0;
    end else begin
      if (11'h557 == _T_12323) begin
        mem_1367 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1368 <= 32'h0;
    end else begin
      if (11'h558 == _T_12323) begin
        mem_1368 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1369 <= 32'h0;
    end else begin
      if (11'h559 == _T_12323) begin
        mem_1369 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1370 <= 32'h0;
    end else begin
      if (11'h55a == _T_12323) begin
        mem_1370 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1371 <= 32'h0;
    end else begin
      if (11'h55b == _T_12323) begin
        mem_1371 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1372 <= 32'h0;
    end else begin
      if (11'h55c == _T_12323) begin
        mem_1372 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1373 <= 32'h0;
    end else begin
      if (11'h55d == _T_12323) begin
        mem_1373 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1374 <= 32'h0;
    end else begin
      if (11'h55e == _T_12323) begin
        mem_1374 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1375 <= 32'h0;
    end else begin
      if (11'h55f == _T_12323) begin
        mem_1375 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1376 <= 32'h0;
    end else begin
      if (11'h560 == _T_12323) begin
        mem_1376 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1377 <= 32'h0;
    end else begin
      if (11'h561 == _T_12323) begin
        mem_1377 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1378 <= 32'h0;
    end else begin
      if (11'h562 == _T_12323) begin
        mem_1378 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1379 <= 32'h0;
    end else begin
      if (11'h563 == _T_12323) begin
        mem_1379 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1380 <= 32'h0;
    end else begin
      if (11'h564 == _T_12323) begin
        mem_1380 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1381 <= 32'h0;
    end else begin
      if (11'h565 == _T_12323) begin
        mem_1381 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1382 <= 32'h0;
    end else begin
      if (11'h566 == _T_12323) begin
        mem_1382 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1383 <= 32'h0;
    end else begin
      if (11'h567 == _T_12323) begin
        mem_1383 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1384 <= 32'h0;
    end else begin
      if (11'h568 == _T_12323) begin
        mem_1384 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1385 <= 32'h0;
    end else begin
      if (11'h569 == _T_12323) begin
        mem_1385 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1386 <= 32'h0;
    end else begin
      if (11'h56a == _T_12323) begin
        mem_1386 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1387 <= 32'h0;
    end else begin
      if (11'h56b == _T_12323) begin
        mem_1387 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1388 <= 32'h0;
    end else begin
      if (11'h56c == _T_12323) begin
        mem_1388 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1389 <= 32'h0;
    end else begin
      if (11'h56d == _T_12323) begin
        mem_1389 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1390 <= 32'h0;
    end else begin
      if (11'h56e == _T_12323) begin
        mem_1390 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1391 <= 32'h0;
    end else begin
      if (11'h56f == _T_12323) begin
        mem_1391 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1392 <= 32'h0;
    end else begin
      if (11'h570 == _T_12323) begin
        mem_1392 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1393 <= 32'h0;
    end else begin
      if (11'h571 == _T_12323) begin
        mem_1393 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1394 <= 32'h0;
    end else begin
      if (11'h572 == _T_12323) begin
        mem_1394 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1395 <= 32'h0;
    end else begin
      if (11'h573 == _T_12323) begin
        mem_1395 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1396 <= 32'h0;
    end else begin
      if (11'h574 == _T_12323) begin
        mem_1396 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1397 <= 32'h0;
    end else begin
      if (11'h575 == _T_12323) begin
        mem_1397 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1398 <= 32'h0;
    end else begin
      if (11'h576 == _T_12323) begin
        mem_1398 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1399 <= 32'h0;
    end else begin
      if (11'h577 == _T_12323) begin
        mem_1399 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1400 <= 32'h0;
    end else begin
      if (11'h578 == _T_12323) begin
        mem_1400 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1401 <= 32'h0;
    end else begin
      if (11'h579 == _T_12323) begin
        mem_1401 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1402 <= 32'h0;
    end else begin
      if (11'h57a == _T_12323) begin
        mem_1402 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1403 <= 32'h0;
    end else begin
      if (11'h57b == _T_12323) begin
        mem_1403 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1404 <= 32'h0;
    end else begin
      if (11'h57c == _T_12323) begin
        mem_1404 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1405 <= 32'h0;
    end else begin
      if (11'h57d == _T_12323) begin
        mem_1405 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1406 <= 32'h0;
    end else begin
      if (11'h57e == _T_12323) begin
        mem_1406 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1407 <= 32'h0;
    end else begin
      if (11'h57f == _T_12323) begin
        mem_1407 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1408 <= 32'h0;
    end else begin
      if (11'h580 == _T_12323) begin
        mem_1408 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1409 <= 32'h0;
    end else begin
      if (11'h581 == _T_12323) begin
        mem_1409 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1410 <= 32'h0;
    end else begin
      if (11'h582 == _T_12323) begin
        mem_1410 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1411 <= 32'h0;
    end else begin
      if (11'h583 == _T_12323) begin
        mem_1411 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1412 <= 32'h0;
    end else begin
      if (11'h584 == _T_12323) begin
        mem_1412 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1413 <= 32'h0;
    end else begin
      if (11'h585 == _T_12323) begin
        mem_1413 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1414 <= 32'h0;
    end else begin
      if (11'h586 == _T_12323) begin
        mem_1414 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1415 <= 32'h0;
    end else begin
      if (11'h587 == _T_12323) begin
        mem_1415 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1416 <= 32'h0;
    end else begin
      if (11'h588 == _T_12323) begin
        mem_1416 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1417 <= 32'h0;
    end else begin
      if (11'h589 == _T_12323) begin
        mem_1417 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1418 <= 32'h0;
    end else begin
      if (11'h58a == _T_12323) begin
        mem_1418 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1419 <= 32'h0;
    end else begin
      if (11'h58b == _T_12323) begin
        mem_1419 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1420 <= 32'h0;
    end else begin
      if (11'h58c == _T_12323) begin
        mem_1420 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1421 <= 32'h0;
    end else begin
      if (11'h58d == _T_12323) begin
        mem_1421 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1422 <= 32'h0;
    end else begin
      if (11'h58e == _T_12323) begin
        mem_1422 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1423 <= 32'h0;
    end else begin
      if (11'h58f == _T_12323) begin
        mem_1423 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1424 <= 32'h0;
    end else begin
      if (11'h590 == _T_12323) begin
        mem_1424 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1425 <= 32'h0;
    end else begin
      if (11'h591 == _T_12323) begin
        mem_1425 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1426 <= 32'h0;
    end else begin
      if (11'h592 == _T_12323) begin
        mem_1426 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1427 <= 32'h0;
    end else begin
      if (11'h593 == _T_12323) begin
        mem_1427 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1428 <= 32'h0;
    end else begin
      if (11'h594 == _T_12323) begin
        mem_1428 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1429 <= 32'h0;
    end else begin
      if (11'h595 == _T_12323) begin
        mem_1429 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1430 <= 32'h0;
    end else begin
      if (11'h596 == _T_12323) begin
        mem_1430 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1431 <= 32'h0;
    end else begin
      if (11'h597 == _T_12323) begin
        mem_1431 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1432 <= 32'h0;
    end else begin
      if (11'h598 == _T_12323) begin
        mem_1432 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1433 <= 32'h0;
    end else begin
      if (11'h599 == _T_12323) begin
        mem_1433 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1434 <= 32'h0;
    end else begin
      if (11'h59a == _T_12323) begin
        mem_1434 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1435 <= 32'h0;
    end else begin
      if (11'h59b == _T_12323) begin
        mem_1435 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1436 <= 32'h0;
    end else begin
      if (11'h59c == _T_12323) begin
        mem_1436 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1437 <= 32'h0;
    end else begin
      if (11'h59d == _T_12323) begin
        mem_1437 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1438 <= 32'h0;
    end else begin
      if (11'h59e == _T_12323) begin
        mem_1438 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1439 <= 32'h0;
    end else begin
      if (11'h59f == _T_12323) begin
        mem_1439 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1440 <= 32'h0;
    end else begin
      if (11'h5a0 == _T_12323) begin
        mem_1440 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1441 <= 32'h0;
    end else begin
      if (11'h5a1 == _T_12323) begin
        mem_1441 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1442 <= 32'h0;
    end else begin
      if (11'h5a2 == _T_12323) begin
        mem_1442 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1443 <= 32'h0;
    end else begin
      if (11'h5a3 == _T_12323) begin
        mem_1443 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1444 <= 32'h0;
    end else begin
      if (11'h5a4 == _T_12323) begin
        mem_1444 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1445 <= 32'h0;
    end else begin
      if (11'h5a5 == _T_12323) begin
        mem_1445 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1446 <= 32'h0;
    end else begin
      if (11'h5a6 == _T_12323) begin
        mem_1446 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1447 <= 32'h0;
    end else begin
      if (11'h5a7 == _T_12323) begin
        mem_1447 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1448 <= 32'h0;
    end else begin
      if (11'h5a8 == _T_12323) begin
        mem_1448 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1449 <= 32'h0;
    end else begin
      if (11'h5a9 == _T_12323) begin
        mem_1449 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1450 <= 32'h0;
    end else begin
      if (11'h5aa == _T_12323) begin
        mem_1450 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1451 <= 32'h0;
    end else begin
      if (11'h5ab == _T_12323) begin
        mem_1451 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1452 <= 32'h0;
    end else begin
      if (11'h5ac == _T_12323) begin
        mem_1452 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1453 <= 32'h0;
    end else begin
      if (11'h5ad == _T_12323) begin
        mem_1453 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1454 <= 32'h0;
    end else begin
      if (11'h5ae == _T_12323) begin
        mem_1454 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1455 <= 32'h0;
    end else begin
      if (11'h5af == _T_12323) begin
        mem_1455 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1456 <= 32'h0;
    end else begin
      if (11'h5b0 == _T_12323) begin
        mem_1456 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1457 <= 32'h0;
    end else begin
      if (11'h5b1 == _T_12323) begin
        mem_1457 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1458 <= 32'h0;
    end else begin
      if (11'h5b2 == _T_12323) begin
        mem_1458 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1459 <= 32'h0;
    end else begin
      if (11'h5b3 == _T_12323) begin
        mem_1459 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1460 <= 32'h0;
    end else begin
      if (11'h5b4 == _T_12323) begin
        mem_1460 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1461 <= 32'h0;
    end else begin
      if (11'h5b5 == _T_12323) begin
        mem_1461 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1462 <= 32'h0;
    end else begin
      if (11'h5b6 == _T_12323) begin
        mem_1462 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1463 <= 32'h0;
    end else begin
      if (11'h5b7 == _T_12323) begin
        mem_1463 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1464 <= 32'h0;
    end else begin
      if (11'h5b8 == _T_12323) begin
        mem_1464 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1465 <= 32'h0;
    end else begin
      if (11'h5b9 == _T_12323) begin
        mem_1465 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1466 <= 32'h0;
    end else begin
      if (11'h5ba == _T_12323) begin
        mem_1466 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1467 <= 32'h0;
    end else begin
      if (11'h5bb == _T_12323) begin
        mem_1467 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1468 <= 32'h0;
    end else begin
      if (11'h5bc == _T_12323) begin
        mem_1468 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1469 <= 32'h0;
    end else begin
      if (11'h5bd == _T_12323) begin
        mem_1469 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1470 <= 32'h0;
    end else begin
      if (11'h5be == _T_12323) begin
        mem_1470 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1471 <= 32'h0;
    end else begin
      if (11'h5bf == _T_12323) begin
        mem_1471 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1472 <= 32'h0;
    end else begin
      if (11'h5c0 == _T_12323) begin
        mem_1472 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1473 <= 32'h0;
    end else begin
      if (11'h5c1 == _T_12323) begin
        mem_1473 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1474 <= 32'h0;
    end else begin
      if (11'h5c2 == _T_12323) begin
        mem_1474 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1475 <= 32'h0;
    end else begin
      if (11'h5c3 == _T_12323) begin
        mem_1475 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1476 <= 32'h0;
    end else begin
      if (11'h5c4 == _T_12323) begin
        mem_1476 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1477 <= 32'h0;
    end else begin
      if (11'h5c5 == _T_12323) begin
        mem_1477 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1478 <= 32'h0;
    end else begin
      if (11'h5c6 == _T_12323) begin
        mem_1478 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1479 <= 32'h0;
    end else begin
      if (11'h5c7 == _T_12323) begin
        mem_1479 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1480 <= 32'h0;
    end else begin
      if (11'h5c8 == _T_12323) begin
        mem_1480 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1481 <= 32'h0;
    end else begin
      if (11'h5c9 == _T_12323) begin
        mem_1481 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1482 <= 32'h0;
    end else begin
      if (11'h5ca == _T_12323) begin
        mem_1482 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1483 <= 32'h0;
    end else begin
      if (11'h5cb == _T_12323) begin
        mem_1483 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1484 <= 32'h0;
    end else begin
      if (11'h5cc == _T_12323) begin
        mem_1484 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1485 <= 32'h0;
    end else begin
      if (11'h5cd == _T_12323) begin
        mem_1485 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1486 <= 32'h0;
    end else begin
      if (11'h5ce == _T_12323) begin
        mem_1486 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1487 <= 32'h0;
    end else begin
      if (11'h5cf == _T_12323) begin
        mem_1487 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1488 <= 32'h0;
    end else begin
      if (11'h5d0 == _T_12323) begin
        mem_1488 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1489 <= 32'h0;
    end else begin
      if (11'h5d1 == _T_12323) begin
        mem_1489 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1490 <= 32'h0;
    end else begin
      if (11'h5d2 == _T_12323) begin
        mem_1490 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1491 <= 32'h0;
    end else begin
      if (11'h5d3 == _T_12323) begin
        mem_1491 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1492 <= 32'h0;
    end else begin
      if (11'h5d4 == _T_12323) begin
        mem_1492 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1493 <= 32'h0;
    end else begin
      if (11'h5d5 == _T_12323) begin
        mem_1493 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1494 <= 32'h0;
    end else begin
      if (11'h5d6 == _T_12323) begin
        mem_1494 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1495 <= 32'h0;
    end else begin
      if (11'h5d7 == _T_12323) begin
        mem_1495 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1496 <= 32'h0;
    end else begin
      if (11'h5d8 == _T_12323) begin
        mem_1496 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1497 <= 32'h0;
    end else begin
      if (11'h5d9 == _T_12323) begin
        mem_1497 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1498 <= 32'h0;
    end else begin
      if (11'h5da == _T_12323) begin
        mem_1498 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1499 <= 32'h0;
    end else begin
      if (11'h5db == _T_12323) begin
        mem_1499 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1500 <= 32'h0;
    end else begin
      if (11'h5dc == _T_12323) begin
        mem_1500 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1501 <= 32'h0;
    end else begin
      if (11'h5dd == _T_12323) begin
        mem_1501 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1502 <= 32'h0;
    end else begin
      if (11'h5de == _T_12323) begin
        mem_1502 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1503 <= 32'h0;
    end else begin
      if (11'h5df == _T_12323) begin
        mem_1503 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1504 <= 32'h0;
    end else begin
      if (11'h5e0 == _T_12323) begin
        mem_1504 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1505 <= 32'h0;
    end else begin
      if (11'h5e1 == _T_12323) begin
        mem_1505 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1506 <= 32'h0;
    end else begin
      if (11'h5e2 == _T_12323) begin
        mem_1506 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1507 <= 32'h0;
    end else begin
      if (11'h5e3 == _T_12323) begin
        mem_1507 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1508 <= 32'h0;
    end else begin
      if (11'h5e4 == _T_12323) begin
        mem_1508 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1509 <= 32'h0;
    end else begin
      if (11'h5e5 == _T_12323) begin
        mem_1509 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1510 <= 32'h0;
    end else begin
      if (11'h5e6 == _T_12323) begin
        mem_1510 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1511 <= 32'h0;
    end else begin
      if (11'h5e7 == _T_12323) begin
        mem_1511 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1512 <= 32'h0;
    end else begin
      if (11'h5e8 == _T_12323) begin
        mem_1512 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1513 <= 32'h0;
    end else begin
      if (11'h5e9 == _T_12323) begin
        mem_1513 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1514 <= 32'h0;
    end else begin
      if (11'h5ea == _T_12323) begin
        mem_1514 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1515 <= 32'h0;
    end else begin
      if (11'h5eb == _T_12323) begin
        mem_1515 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1516 <= 32'h0;
    end else begin
      if (11'h5ec == _T_12323) begin
        mem_1516 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1517 <= 32'h0;
    end else begin
      if (11'h5ed == _T_12323) begin
        mem_1517 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1518 <= 32'h0;
    end else begin
      if (11'h5ee == _T_12323) begin
        mem_1518 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1519 <= 32'h0;
    end else begin
      if (11'h5ef == _T_12323) begin
        mem_1519 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1520 <= 32'h0;
    end else begin
      if (11'h5f0 == _T_12323) begin
        mem_1520 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1521 <= 32'h0;
    end else begin
      if (11'h5f1 == _T_12323) begin
        mem_1521 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1522 <= 32'h0;
    end else begin
      if (11'h5f2 == _T_12323) begin
        mem_1522 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1523 <= 32'h0;
    end else begin
      if (11'h5f3 == _T_12323) begin
        mem_1523 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1524 <= 32'h0;
    end else begin
      if (11'h5f4 == _T_12323) begin
        mem_1524 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1525 <= 32'h0;
    end else begin
      if (11'h5f5 == _T_12323) begin
        mem_1525 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1526 <= 32'h0;
    end else begin
      if (11'h5f6 == _T_12323) begin
        mem_1526 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1527 <= 32'h0;
    end else begin
      if (11'h5f7 == _T_12323) begin
        mem_1527 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1528 <= 32'h0;
    end else begin
      if (11'h5f8 == _T_12323) begin
        mem_1528 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1529 <= 32'h0;
    end else begin
      if (11'h5f9 == _T_12323) begin
        mem_1529 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1530 <= 32'h0;
    end else begin
      if (11'h5fa == _T_12323) begin
        mem_1530 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1531 <= 32'h0;
    end else begin
      if (11'h5fb == _T_12323) begin
        mem_1531 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1532 <= 32'h0;
    end else begin
      if (11'h5fc == _T_12323) begin
        mem_1532 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1533 <= 32'h0;
    end else begin
      if (11'h5fd == _T_12323) begin
        mem_1533 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1534 <= 32'h0;
    end else begin
      if (11'h5fe == _T_12323) begin
        mem_1534 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1535 <= 32'h0;
    end else begin
      if (11'h5ff == _T_12323) begin
        mem_1535 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1536 <= 32'h0;
    end else begin
      if (11'h600 == _T_12323) begin
        mem_1536 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1537 <= 32'h0;
    end else begin
      if (11'h601 == _T_12323) begin
        mem_1537 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1538 <= 32'h0;
    end else begin
      if (11'h602 == _T_12323) begin
        mem_1538 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1539 <= 32'h0;
    end else begin
      if (11'h603 == _T_12323) begin
        mem_1539 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1540 <= 32'h0;
    end else begin
      if (11'h604 == _T_12323) begin
        mem_1540 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1541 <= 32'h0;
    end else begin
      if (11'h605 == _T_12323) begin
        mem_1541 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1542 <= 32'h0;
    end else begin
      if (11'h606 == _T_12323) begin
        mem_1542 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1543 <= 32'h0;
    end else begin
      if (11'h607 == _T_12323) begin
        mem_1543 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1544 <= 32'h0;
    end else begin
      if (11'h608 == _T_12323) begin
        mem_1544 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1545 <= 32'h0;
    end else begin
      if (11'h609 == _T_12323) begin
        mem_1545 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1546 <= 32'h0;
    end else begin
      if (11'h60a == _T_12323) begin
        mem_1546 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1547 <= 32'h0;
    end else begin
      if (11'h60b == _T_12323) begin
        mem_1547 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1548 <= 32'h0;
    end else begin
      if (11'h60c == _T_12323) begin
        mem_1548 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1549 <= 32'h0;
    end else begin
      if (11'h60d == _T_12323) begin
        mem_1549 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1550 <= 32'h0;
    end else begin
      if (11'h60e == _T_12323) begin
        mem_1550 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1551 <= 32'h0;
    end else begin
      if (11'h60f == _T_12323) begin
        mem_1551 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1552 <= 32'h0;
    end else begin
      if (11'h610 == _T_12323) begin
        mem_1552 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1553 <= 32'h0;
    end else begin
      if (11'h611 == _T_12323) begin
        mem_1553 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1554 <= 32'h0;
    end else begin
      if (11'h612 == _T_12323) begin
        mem_1554 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1555 <= 32'h0;
    end else begin
      if (11'h613 == _T_12323) begin
        mem_1555 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1556 <= 32'h0;
    end else begin
      if (11'h614 == _T_12323) begin
        mem_1556 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1557 <= 32'h0;
    end else begin
      if (11'h615 == _T_12323) begin
        mem_1557 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1558 <= 32'h0;
    end else begin
      if (11'h616 == _T_12323) begin
        mem_1558 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1559 <= 32'h0;
    end else begin
      if (11'h617 == _T_12323) begin
        mem_1559 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1560 <= 32'h0;
    end else begin
      if (11'h618 == _T_12323) begin
        mem_1560 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1561 <= 32'h0;
    end else begin
      if (11'h619 == _T_12323) begin
        mem_1561 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1562 <= 32'h0;
    end else begin
      if (11'h61a == _T_12323) begin
        mem_1562 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1563 <= 32'h0;
    end else begin
      if (11'h61b == _T_12323) begin
        mem_1563 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1564 <= 32'h0;
    end else begin
      if (11'h61c == _T_12323) begin
        mem_1564 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1565 <= 32'h0;
    end else begin
      if (11'h61d == _T_12323) begin
        mem_1565 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1566 <= 32'h0;
    end else begin
      if (11'h61e == _T_12323) begin
        mem_1566 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1567 <= 32'h0;
    end else begin
      if (11'h61f == _T_12323) begin
        mem_1567 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1568 <= 32'h0;
    end else begin
      if (11'h620 == _T_12323) begin
        mem_1568 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1569 <= 32'h0;
    end else begin
      if (11'h621 == _T_12323) begin
        mem_1569 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1570 <= 32'h0;
    end else begin
      if (11'h622 == _T_12323) begin
        mem_1570 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1571 <= 32'h0;
    end else begin
      if (11'h623 == _T_12323) begin
        mem_1571 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1572 <= 32'h0;
    end else begin
      if (11'h624 == _T_12323) begin
        mem_1572 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1573 <= 32'h0;
    end else begin
      if (11'h625 == _T_12323) begin
        mem_1573 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1574 <= 32'h0;
    end else begin
      if (11'h626 == _T_12323) begin
        mem_1574 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1575 <= 32'h0;
    end else begin
      if (11'h627 == _T_12323) begin
        mem_1575 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1576 <= 32'h0;
    end else begin
      if (11'h628 == _T_12323) begin
        mem_1576 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1577 <= 32'h0;
    end else begin
      if (11'h629 == _T_12323) begin
        mem_1577 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1578 <= 32'h0;
    end else begin
      if (11'h62a == _T_12323) begin
        mem_1578 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1579 <= 32'h0;
    end else begin
      if (11'h62b == _T_12323) begin
        mem_1579 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1580 <= 32'h0;
    end else begin
      if (11'h62c == _T_12323) begin
        mem_1580 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1581 <= 32'h0;
    end else begin
      if (11'h62d == _T_12323) begin
        mem_1581 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1582 <= 32'h0;
    end else begin
      if (11'h62e == _T_12323) begin
        mem_1582 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1583 <= 32'h0;
    end else begin
      if (11'h62f == _T_12323) begin
        mem_1583 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1584 <= 32'h0;
    end else begin
      if (11'h630 == _T_12323) begin
        mem_1584 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1585 <= 32'h0;
    end else begin
      if (11'h631 == _T_12323) begin
        mem_1585 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1586 <= 32'h0;
    end else begin
      if (11'h632 == _T_12323) begin
        mem_1586 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1587 <= 32'h0;
    end else begin
      if (11'h633 == _T_12323) begin
        mem_1587 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1588 <= 32'h0;
    end else begin
      if (11'h634 == _T_12323) begin
        mem_1588 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1589 <= 32'h0;
    end else begin
      if (11'h635 == _T_12323) begin
        mem_1589 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1590 <= 32'h0;
    end else begin
      if (11'h636 == _T_12323) begin
        mem_1590 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1591 <= 32'h0;
    end else begin
      if (11'h637 == _T_12323) begin
        mem_1591 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1592 <= 32'h0;
    end else begin
      if (11'h638 == _T_12323) begin
        mem_1592 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1593 <= 32'h0;
    end else begin
      if (11'h639 == _T_12323) begin
        mem_1593 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1594 <= 32'h0;
    end else begin
      if (11'h63a == _T_12323) begin
        mem_1594 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1595 <= 32'h0;
    end else begin
      if (11'h63b == _T_12323) begin
        mem_1595 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1596 <= 32'h0;
    end else begin
      if (11'h63c == _T_12323) begin
        mem_1596 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1597 <= 32'h0;
    end else begin
      if (11'h63d == _T_12323) begin
        mem_1597 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1598 <= 32'h0;
    end else begin
      if (11'h63e == _T_12323) begin
        mem_1598 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1599 <= 32'h0;
    end else begin
      if (11'h63f == _T_12323) begin
        mem_1599 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1600 <= 32'h0;
    end else begin
      if (11'h640 == _T_12323) begin
        mem_1600 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1601 <= 32'h0;
    end else begin
      if (11'h641 == _T_12323) begin
        mem_1601 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1602 <= 32'h0;
    end else begin
      if (11'h642 == _T_12323) begin
        mem_1602 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1603 <= 32'h0;
    end else begin
      if (11'h643 == _T_12323) begin
        mem_1603 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1604 <= 32'h0;
    end else begin
      if (11'h644 == _T_12323) begin
        mem_1604 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1605 <= 32'h0;
    end else begin
      if (11'h645 == _T_12323) begin
        mem_1605 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1606 <= 32'h0;
    end else begin
      if (11'h646 == _T_12323) begin
        mem_1606 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1607 <= 32'h0;
    end else begin
      if (11'h647 == _T_12323) begin
        mem_1607 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1608 <= 32'h0;
    end else begin
      if (11'h648 == _T_12323) begin
        mem_1608 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1609 <= 32'h0;
    end else begin
      if (11'h649 == _T_12323) begin
        mem_1609 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1610 <= 32'h0;
    end else begin
      if (11'h64a == _T_12323) begin
        mem_1610 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1611 <= 32'h0;
    end else begin
      if (11'h64b == _T_12323) begin
        mem_1611 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1612 <= 32'h0;
    end else begin
      if (11'h64c == _T_12323) begin
        mem_1612 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1613 <= 32'h0;
    end else begin
      if (11'h64d == _T_12323) begin
        mem_1613 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1614 <= 32'h0;
    end else begin
      if (11'h64e == _T_12323) begin
        mem_1614 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1615 <= 32'h0;
    end else begin
      if (11'h64f == _T_12323) begin
        mem_1615 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1616 <= 32'h0;
    end else begin
      if (11'h650 == _T_12323) begin
        mem_1616 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1617 <= 32'h0;
    end else begin
      if (11'h651 == _T_12323) begin
        mem_1617 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1618 <= 32'h0;
    end else begin
      if (11'h652 == _T_12323) begin
        mem_1618 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1619 <= 32'h0;
    end else begin
      if (11'h653 == _T_12323) begin
        mem_1619 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1620 <= 32'h0;
    end else begin
      if (11'h654 == _T_12323) begin
        mem_1620 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1621 <= 32'h0;
    end else begin
      if (11'h655 == _T_12323) begin
        mem_1621 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1622 <= 32'h0;
    end else begin
      if (11'h656 == _T_12323) begin
        mem_1622 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1623 <= 32'h0;
    end else begin
      if (11'h657 == _T_12323) begin
        mem_1623 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1624 <= 32'h0;
    end else begin
      if (11'h658 == _T_12323) begin
        mem_1624 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1625 <= 32'h0;
    end else begin
      if (11'h659 == _T_12323) begin
        mem_1625 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1626 <= 32'h0;
    end else begin
      if (11'h65a == _T_12323) begin
        mem_1626 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1627 <= 32'h0;
    end else begin
      if (11'h65b == _T_12323) begin
        mem_1627 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1628 <= 32'h0;
    end else begin
      if (11'h65c == _T_12323) begin
        mem_1628 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1629 <= 32'h0;
    end else begin
      if (11'h65d == _T_12323) begin
        mem_1629 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1630 <= 32'h0;
    end else begin
      if (11'h65e == _T_12323) begin
        mem_1630 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1631 <= 32'h0;
    end else begin
      if (11'h65f == _T_12323) begin
        mem_1631 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1632 <= 32'h0;
    end else begin
      if (11'h660 == _T_12323) begin
        mem_1632 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1633 <= 32'h0;
    end else begin
      if (11'h661 == _T_12323) begin
        mem_1633 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1634 <= 32'h0;
    end else begin
      if (11'h662 == _T_12323) begin
        mem_1634 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1635 <= 32'h0;
    end else begin
      if (11'h663 == _T_12323) begin
        mem_1635 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1636 <= 32'h0;
    end else begin
      if (11'h664 == _T_12323) begin
        mem_1636 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1637 <= 32'h0;
    end else begin
      if (11'h665 == _T_12323) begin
        mem_1637 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1638 <= 32'h0;
    end else begin
      if (11'h666 == _T_12323) begin
        mem_1638 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1639 <= 32'h0;
    end else begin
      if (11'h667 == _T_12323) begin
        mem_1639 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1640 <= 32'h0;
    end else begin
      if (11'h668 == _T_12323) begin
        mem_1640 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1641 <= 32'h0;
    end else begin
      if (11'h669 == _T_12323) begin
        mem_1641 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1642 <= 32'h0;
    end else begin
      if (11'h66a == _T_12323) begin
        mem_1642 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1643 <= 32'h0;
    end else begin
      if (11'h66b == _T_12323) begin
        mem_1643 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1644 <= 32'h0;
    end else begin
      if (11'h66c == _T_12323) begin
        mem_1644 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1645 <= 32'h0;
    end else begin
      if (11'h66d == _T_12323) begin
        mem_1645 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1646 <= 32'h0;
    end else begin
      if (11'h66e == _T_12323) begin
        mem_1646 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1647 <= 32'h0;
    end else begin
      if (11'h66f == _T_12323) begin
        mem_1647 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1648 <= 32'h0;
    end else begin
      if (11'h670 == _T_12323) begin
        mem_1648 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1649 <= 32'h0;
    end else begin
      if (11'h671 == _T_12323) begin
        mem_1649 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1650 <= 32'h0;
    end else begin
      if (11'h672 == _T_12323) begin
        mem_1650 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1651 <= 32'h0;
    end else begin
      if (11'h673 == _T_12323) begin
        mem_1651 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1652 <= 32'h0;
    end else begin
      if (11'h674 == _T_12323) begin
        mem_1652 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1653 <= 32'h0;
    end else begin
      if (11'h675 == _T_12323) begin
        mem_1653 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1654 <= 32'h0;
    end else begin
      if (11'h676 == _T_12323) begin
        mem_1654 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1655 <= 32'h0;
    end else begin
      if (11'h677 == _T_12323) begin
        mem_1655 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1656 <= 32'h0;
    end else begin
      if (11'h678 == _T_12323) begin
        mem_1656 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1657 <= 32'h0;
    end else begin
      if (11'h679 == _T_12323) begin
        mem_1657 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1658 <= 32'h0;
    end else begin
      if (11'h67a == _T_12323) begin
        mem_1658 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1659 <= 32'h0;
    end else begin
      if (11'h67b == _T_12323) begin
        mem_1659 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1660 <= 32'h0;
    end else begin
      if (11'h67c == _T_12323) begin
        mem_1660 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1661 <= 32'h0;
    end else begin
      if (11'h67d == _T_12323) begin
        mem_1661 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1662 <= 32'h0;
    end else begin
      if (11'h67e == _T_12323) begin
        mem_1662 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1663 <= 32'h0;
    end else begin
      if (11'h67f == _T_12323) begin
        mem_1663 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1664 <= 32'h0;
    end else begin
      if (11'h680 == _T_12323) begin
        mem_1664 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1665 <= 32'h0;
    end else begin
      if (11'h681 == _T_12323) begin
        mem_1665 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1666 <= 32'h0;
    end else begin
      if (11'h682 == _T_12323) begin
        mem_1666 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1667 <= 32'h0;
    end else begin
      if (11'h683 == _T_12323) begin
        mem_1667 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1668 <= 32'h0;
    end else begin
      if (11'h684 == _T_12323) begin
        mem_1668 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1669 <= 32'h0;
    end else begin
      if (11'h685 == _T_12323) begin
        mem_1669 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1670 <= 32'h0;
    end else begin
      if (11'h686 == _T_12323) begin
        mem_1670 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1671 <= 32'h0;
    end else begin
      if (11'h687 == _T_12323) begin
        mem_1671 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1672 <= 32'h0;
    end else begin
      if (11'h688 == _T_12323) begin
        mem_1672 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1673 <= 32'h0;
    end else begin
      if (11'h689 == _T_12323) begin
        mem_1673 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1674 <= 32'h0;
    end else begin
      if (11'h68a == _T_12323) begin
        mem_1674 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1675 <= 32'h0;
    end else begin
      if (11'h68b == _T_12323) begin
        mem_1675 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1676 <= 32'h0;
    end else begin
      if (11'h68c == _T_12323) begin
        mem_1676 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1677 <= 32'h0;
    end else begin
      if (11'h68d == _T_12323) begin
        mem_1677 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1678 <= 32'h0;
    end else begin
      if (11'h68e == _T_12323) begin
        mem_1678 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1679 <= 32'h0;
    end else begin
      if (11'h68f == _T_12323) begin
        mem_1679 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1680 <= 32'h0;
    end else begin
      if (11'h690 == _T_12323) begin
        mem_1680 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1681 <= 32'h0;
    end else begin
      if (11'h691 == _T_12323) begin
        mem_1681 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1682 <= 32'h0;
    end else begin
      if (11'h692 == _T_12323) begin
        mem_1682 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1683 <= 32'h0;
    end else begin
      if (11'h693 == _T_12323) begin
        mem_1683 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1684 <= 32'h0;
    end else begin
      if (11'h694 == _T_12323) begin
        mem_1684 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1685 <= 32'h0;
    end else begin
      if (11'h695 == _T_12323) begin
        mem_1685 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1686 <= 32'h0;
    end else begin
      if (11'h696 == _T_12323) begin
        mem_1686 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1687 <= 32'h0;
    end else begin
      if (11'h697 == _T_12323) begin
        mem_1687 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1688 <= 32'h0;
    end else begin
      if (11'h698 == _T_12323) begin
        mem_1688 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1689 <= 32'h0;
    end else begin
      if (11'h699 == _T_12323) begin
        mem_1689 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1690 <= 32'h0;
    end else begin
      if (11'h69a == _T_12323) begin
        mem_1690 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1691 <= 32'h0;
    end else begin
      if (11'h69b == _T_12323) begin
        mem_1691 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1692 <= 32'h0;
    end else begin
      if (11'h69c == _T_12323) begin
        mem_1692 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1693 <= 32'h0;
    end else begin
      if (11'h69d == _T_12323) begin
        mem_1693 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1694 <= 32'h0;
    end else begin
      if (11'h69e == _T_12323) begin
        mem_1694 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1695 <= 32'h0;
    end else begin
      if (11'h69f == _T_12323) begin
        mem_1695 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1696 <= 32'h0;
    end else begin
      if (11'h6a0 == _T_12323) begin
        mem_1696 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1697 <= 32'h0;
    end else begin
      if (11'h6a1 == _T_12323) begin
        mem_1697 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1698 <= 32'h0;
    end else begin
      if (11'h6a2 == _T_12323) begin
        mem_1698 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1699 <= 32'h0;
    end else begin
      if (11'h6a3 == _T_12323) begin
        mem_1699 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1700 <= 32'h0;
    end else begin
      if (11'h6a4 == _T_12323) begin
        mem_1700 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1701 <= 32'h0;
    end else begin
      if (11'h6a5 == _T_12323) begin
        mem_1701 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1702 <= 32'h0;
    end else begin
      if (11'h6a6 == _T_12323) begin
        mem_1702 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1703 <= 32'h0;
    end else begin
      if (11'h6a7 == _T_12323) begin
        mem_1703 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1704 <= 32'h0;
    end else begin
      if (11'h6a8 == _T_12323) begin
        mem_1704 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1705 <= 32'h0;
    end else begin
      if (11'h6a9 == _T_12323) begin
        mem_1705 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1706 <= 32'h0;
    end else begin
      if (11'h6aa == _T_12323) begin
        mem_1706 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1707 <= 32'h0;
    end else begin
      if (11'h6ab == _T_12323) begin
        mem_1707 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1708 <= 32'h0;
    end else begin
      if (11'h6ac == _T_12323) begin
        mem_1708 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1709 <= 32'h0;
    end else begin
      if (11'h6ad == _T_12323) begin
        mem_1709 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1710 <= 32'h0;
    end else begin
      if (11'h6ae == _T_12323) begin
        mem_1710 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1711 <= 32'h0;
    end else begin
      if (11'h6af == _T_12323) begin
        mem_1711 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1712 <= 32'h0;
    end else begin
      if (11'h6b0 == _T_12323) begin
        mem_1712 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1713 <= 32'h0;
    end else begin
      if (11'h6b1 == _T_12323) begin
        mem_1713 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1714 <= 32'h0;
    end else begin
      if (11'h6b2 == _T_12323) begin
        mem_1714 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1715 <= 32'h0;
    end else begin
      if (11'h6b3 == _T_12323) begin
        mem_1715 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1716 <= 32'h0;
    end else begin
      if (11'h6b4 == _T_12323) begin
        mem_1716 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1717 <= 32'h0;
    end else begin
      if (11'h6b5 == _T_12323) begin
        mem_1717 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1718 <= 32'h0;
    end else begin
      if (11'h6b6 == _T_12323) begin
        mem_1718 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1719 <= 32'h0;
    end else begin
      if (11'h6b7 == _T_12323) begin
        mem_1719 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1720 <= 32'h0;
    end else begin
      if (11'h6b8 == _T_12323) begin
        mem_1720 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1721 <= 32'h0;
    end else begin
      if (11'h6b9 == _T_12323) begin
        mem_1721 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1722 <= 32'h0;
    end else begin
      if (11'h6ba == _T_12323) begin
        mem_1722 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1723 <= 32'h0;
    end else begin
      if (11'h6bb == _T_12323) begin
        mem_1723 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1724 <= 32'h0;
    end else begin
      if (11'h6bc == _T_12323) begin
        mem_1724 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1725 <= 32'h0;
    end else begin
      if (11'h6bd == _T_12323) begin
        mem_1725 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1726 <= 32'h0;
    end else begin
      if (11'h6be == _T_12323) begin
        mem_1726 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1727 <= 32'h0;
    end else begin
      if (11'h6bf == _T_12323) begin
        mem_1727 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1728 <= 32'h0;
    end else begin
      if (11'h6c0 == _T_12323) begin
        mem_1728 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1729 <= 32'h0;
    end else begin
      if (11'h6c1 == _T_12323) begin
        mem_1729 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1730 <= 32'h0;
    end else begin
      if (11'h6c2 == _T_12323) begin
        mem_1730 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1731 <= 32'h0;
    end else begin
      if (11'h6c3 == _T_12323) begin
        mem_1731 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1732 <= 32'h0;
    end else begin
      if (11'h6c4 == _T_12323) begin
        mem_1732 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1733 <= 32'h0;
    end else begin
      if (11'h6c5 == _T_12323) begin
        mem_1733 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1734 <= 32'h0;
    end else begin
      if (11'h6c6 == _T_12323) begin
        mem_1734 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1735 <= 32'h0;
    end else begin
      if (11'h6c7 == _T_12323) begin
        mem_1735 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1736 <= 32'h0;
    end else begin
      if (11'h6c8 == _T_12323) begin
        mem_1736 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1737 <= 32'h0;
    end else begin
      if (11'h6c9 == _T_12323) begin
        mem_1737 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1738 <= 32'h0;
    end else begin
      if (11'h6ca == _T_12323) begin
        mem_1738 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1739 <= 32'h0;
    end else begin
      if (11'h6cb == _T_12323) begin
        mem_1739 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1740 <= 32'h0;
    end else begin
      if (11'h6cc == _T_12323) begin
        mem_1740 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1741 <= 32'h0;
    end else begin
      if (11'h6cd == _T_12323) begin
        mem_1741 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1742 <= 32'h0;
    end else begin
      if (11'h6ce == _T_12323) begin
        mem_1742 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1743 <= 32'h0;
    end else begin
      if (11'h6cf == _T_12323) begin
        mem_1743 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1744 <= 32'h0;
    end else begin
      if (11'h6d0 == _T_12323) begin
        mem_1744 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1745 <= 32'h0;
    end else begin
      if (11'h6d1 == _T_12323) begin
        mem_1745 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1746 <= 32'h0;
    end else begin
      if (11'h6d2 == _T_12323) begin
        mem_1746 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1747 <= 32'h0;
    end else begin
      if (11'h6d3 == _T_12323) begin
        mem_1747 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1748 <= 32'h0;
    end else begin
      if (11'h6d4 == _T_12323) begin
        mem_1748 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1749 <= 32'h0;
    end else begin
      if (11'h6d5 == _T_12323) begin
        mem_1749 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1750 <= 32'h0;
    end else begin
      if (11'h6d6 == _T_12323) begin
        mem_1750 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1751 <= 32'h0;
    end else begin
      if (11'h6d7 == _T_12323) begin
        mem_1751 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1752 <= 32'h0;
    end else begin
      if (11'h6d8 == _T_12323) begin
        mem_1752 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1753 <= 32'h0;
    end else begin
      if (11'h6d9 == _T_12323) begin
        mem_1753 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1754 <= 32'h0;
    end else begin
      if (11'h6da == _T_12323) begin
        mem_1754 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1755 <= 32'h0;
    end else begin
      if (11'h6db == _T_12323) begin
        mem_1755 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1756 <= 32'h0;
    end else begin
      if (11'h6dc == _T_12323) begin
        mem_1756 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1757 <= 32'h0;
    end else begin
      if (11'h6dd == _T_12323) begin
        mem_1757 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1758 <= 32'h0;
    end else begin
      if (11'h6de == _T_12323) begin
        mem_1758 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1759 <= 32'h0;
    end else begin
      if (11'h6df == _T_12323) begin
        mem_1759 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1760 <= 32'h0;
    end else begin
      if (11'h6e0 == _T_12323) begin
        mem_1760 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1761 <= 32'h0;
    end else begin
      if (11'h6e1 == _T_12323) begin
        mem_1761 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1762 <= 32'h0;
    end else begin
      if (11'h6e2 == _T_12323) begin
        mem_1762 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1763 <= 32'h0;
    end else begin
      if (11'h6e3 == _T_12323) begin
        mem_1763 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1764 <= 32'h0;
    end else begin
      if (11'h6e4 == _T_12323) begin
        mem_1764 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1765 <= 32'h0;
    end else begin
      if (11'h6e5 == _T_12323) begin
        mem_1765 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1766 <= 32'h0;
    end else begin
      if (11'h6e6 == _T_12323) begin
        mem_1766 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1767 <= 32'h0;
    end else begin
      if (11'h6e7 == _T_12323) begin
        mem_1767 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1768 <= 32'h0;
    end else begin
      if (11'h6e8 == _T_12323) begin
        mem_1768 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1769 <= 32'h0;
    end else begin
      if (11'h6e9 == _T_12323) begin
        mem_1769 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1770 <= 32'h0;
    end else begin
      if (11'h6ea == _T_12323) begin
        mem_1770 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1771 <= 32'h0;
    end else begin
      if (11'h6eb == _T_12323) begin
        mem_1771 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1772 <= 32'h0;
    end else begin
      if (11'h6ec == _T_12323) begin
        mem_1772 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1773 <= 32'h0;
    end else begin
      if (11'h6ed == _T_12323) begin
        mem_1773 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1774 <= 32'h0;
    end else begin
      if (11'h6ee == _T_12323) begin
        mem_1774 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1775 <= 32'h0;
    end else begin
      if (11'h6ef == _T_12323) begin
        mem_1775 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1776 <= 32'h0;
    end else begin
      if (11'h6f0 == _T_12323) begin
        mem_1776 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1777 <= 32'h0;
    end else begin
      if (11'h6f1 == _T_12323) begin
        mem_1777 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1778 <= 32'h0;
    end else begin
      if (11'h6f2 == _T_12323) begin
        mem_1778 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1779 <= 32'h0;
    end else begin
      if (11'h6f3 == _T_12323) begin
        mem_1779 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1780 <= 32'h0;
    end else begin
      if (11'h6f4 == _T_12323) begin
        mem_1780 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1781 <= 32'h0;
    end else begin
      if (11'h6f5 == _T_12323) begin
        mem_1781 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1782 <= 32'h0;
    end else begin
      if (11'h6f6 == _T_12323) begin
        mem_1782 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1783 <= 32'h0;
    end else begin
      if (11'h6f7 == _T_12323) begin
        mem_1783 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1784 <= 32'h0;
    end else begin
      if (11'h6f8 == _T_12323) begin
        mem_1784 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1785 <= 32'h0;
    end else begin
      if (11'h6f9 == _T_12323) begin
        mem_1785 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1786 <= 32'h0;
    end else begin
      if (11'h6fa == _T_12323) begin
        mem_1786 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1787 <= 32'h0;
    end else begin
      if (11'h6fb == _T_12323) begin
        mem_1787 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1788 <= 32'h0;
    end else begin
      if (11'h6fc == _T_12323) begin
        mem_1788 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1789 <= 32'h0;
    end else begin
      if (11'h6fd == _T_12323) begin
        mem_1789 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1790 <= 32'h0;
    end else begin
      if (11'h6fe == _T_12323) begin
        mem_1790 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1791 <= 32'h0;
    end else begin
      if (11'h6ff == _T_12323) begin
        mem_1791 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1792 <= 32'h0;
    end else begin
      if (11'h700 == _T_12323) begin
        mem_1792 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1793 <= 32'h0;
    end else begin
      if (11'h701 == _T_12323) begin
        mem_1793 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1794 <= 32'h0;
    end else begin
      if (11'h702 == _T_12323) begin
        mem_1794 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1795 <= 32'h0;
    end else begin
      if (11'h703 == _T_12323) begin
        mem_1795 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1796 <= 32'h0;
    end else begin
      if (11'h704 == _T_12323) begin
        mem_1796 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1797 <= 32'h0;
    end else begin
      if (11'h705 == _T_12323) begin
        mem_1797 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1798 <= 32'h0;
    end else begin
      if (11'h706 == _T_12323) begin
        mem_1798 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1799 <= 32'h0;
    end else begin
      if (11'h707 == _T_12323) begin
        mem_1799 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1800 <= 32'h0;
    end else begin
      if (11'h708 == _T_12323) begin
        mem_1800 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1801 <= 32'h0;
    end else begin
      if (11'h709 == _T_12323) begin
        mem_1801 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1802 <= 32'h0;
    end else begin
      if (11'h70a == _T_12323) begin
        mem_1802 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1803 <= 32'h0;
    end else begin
      if (11'h70b == _T_12323) begin
        mem_1803 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1804 <= 32'h0;
    end else begin
      if (11'h70c == _T_12323) begin
        mem_1804 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1805 <= 32'h0;
    end else begin
      if (11'h70d == _T_12323) begin
        mem_1805 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1806 <= 32'h0;
    end else begin
      if (11'h70e == _T_12323) begin
        mem_1806 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1807 <= 32'h0;
    end else begin
      if (11'h70f == _T_12323) begin
        mem_1807 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1808 <= 32'h0;
    end else begin
      if (11'h710 == _T_12323) begin
        mem_1808 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1809 <= 32'h0;
    end else begin
      if (11'h711 == _T_12323) begin
        mem_1809 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1810 <= 32'h0;
    end else begin
      if (11'h712 == _T_12323) begin
        mem_1810 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1811 <= 32'h0;
    end else begin
      if (11'h713 == _T_12323) begin
        mem_1811 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1812 <= 32'h0;
    end else begin
      if (11'h714 == _T_12323) begin
        mem_1812 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1813 <= 32'h0;
    end else begin
      if (11'h715 == _T_12323) begin
        mem_1813 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1814 <= 32'h0;
    end else begin
      if (11'h716 == _T_12323) begin
        mem_1814 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1815 <= 32'h0;
    end else begin
      if (11'h717 == _T_12323) begin
        mem_1815 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1816 <= 32'h0;
    end else begin
      if (11'h718 == _T_12323) begin
        mem_1816 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1817 <= 32'h0;
    end else begin
      if (11'h719 == _T_12323) begin
        mem_1817 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1818 <= 32'h0;
    end else begin
      if (11'h71a == _T_12323) begin
        mem_1818 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1819 <= 32'h0;
    end else begin
      if (11'h71b == _T_12323) begin
        mem_1819 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1820 <= 32'h0;
    end else begin
      if (11'h71c == _T_12323) begin
        mem_1820 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1821 <= 32'h0;
    end else begin
      if (11'h71d == _T_12323) begin
        mem_1821 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1822 <= 32'h0;
    end else begin
      if (11'h71e == _T_12323) begin
        mem_1822 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1823 <= 32'h0;
    end else begin
      if (11'h71f == _T_12323) begin
        mem_1823 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1824 <= 32'h0;
    end else begin
      if (11'h720 == _T_12323) begin
        mem_1824 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1825 <= 32'h0;
    end else begin
      if (11'h721 == _T_12323) begin
        mem_1825 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1826 <= 32'h0;
    end else begin
      if (11'h722 == _T_12323) begin
        mem_1826 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1827 <= 32'h0;
    end else begin
      if (11'h723 == _T_12323) begin
        mem_1827 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1828 <= 32'h0;
    end else begin
      if (11'h724 == _T_12323) begin
        mem_1828 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1829 <= 32'h0;
    end else begin
      if (11'h725 == _T_12323) begin
        mem_1829 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1830 <= 32'h0;
    end else begin
      if (11'h726 == _T_12323) begin
        mem_1830 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1831 <= 32'h0;
    end else begin
      if (11'h727 == _T_12323) begin
        mem_1831 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1832 <= 32'h0;
    end else begin
      if (11'h728 == _T_12323) begin
        mem_1832 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1833 <= 32'h0;
    end else begin
      if (11'h729 == _T_12323) begin
        mem_1833 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1834 <= 32'h0;
    end else begin
      if (11'h72a == _T_12323) begin
        mem_1834 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1835 <= 32'h0;
    end else begin
      if (11'h72b == _T_12323) begin
        mem_1835 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1836 <= 32'h0;
    end else begin
      if (11'h72c == _T_12323) begin
        mem_1836 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1837 <= 32'h0;
    end else begin
      if (11'h72d == _T_12323) begin
        mem_1837 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1838 <= 32'h0;
    end else begin
      if (11'h72e == _T_12323) begin
        mem_1838 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1839 <= 32'h0;
    end else begin
      if (11'h72f == _T_12323) begin
        mem_1839 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1840 <= 32'h0;
    end else begin
      if (11'h730 == _T_12323) begin
        mem_1840 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1841 <= 32'h0;
    end else begin
      if (11'h731 == _T_12323) begin
        mem_1841 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1842 <= 32'h0;
    end else begin
      if (11'h732 == _T_12323) begin
        mem_1842 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1843 <= 32'h0;
    end else begin
      if (11'h733 == _T_12323) begin
        mem_1843 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1844 <= 32'h0;
    end else begin
      if (11'h734 == _T_12323) begin
        mem_1844 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1845 <= 32'h0;
    end else begin
      if (11'h735 == _T_12323) begin
        mem_1845 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1846 <= 32'h0;
    end else begin
      if (11'h736 == _T_12323) begin
        mem_1846 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1847 <= 32'h0;
    end else begin
      if (11'h737 == _T_12323) begin
        mem_1847 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1848 <= 32'h0;
    end else begin
      if (11'h738 == _T_12323) begin
        mem_1848 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1849 <= 32'h0;
    end else begin
      if (11'h739 == _T_12323) begin
        mem_1849 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1850 <= 32'h0;
    end else begin
      if (11'h73a == _T_12323) begin
        mem_1850 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1851 <= 32'h0;
    end else begin
      if (11'h73b == _T_12323) begin
        mem_1851 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1852 <= 32'h0;
    end else begin
      if (11'h73c == _T_12323) begin
        mem_1852 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1853 <= 32'h0;
    end else begin
      if (11'h73d == _T_12323) begin
        mem_1853 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1854 <= 32'h0;
    end else begin
      if (11'h73e == _T_12323) begin
        mem_1854 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1855 <= 32'h0;
    end else begin
      if (11'h73f == _T_12323) begin
        mem_1855 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1856 <= 32'h0;
    end else begin
      if (11'h740 == _T_12323) begin
        mem_1856 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1857 <= 32'h0;
    end else begin
      if (11'h741 == _T_12323) begin
        mem_1857 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1858 <= 32'h0;
    end else begin
      if (11'h742 == _T_12323) begin
        mem_1858 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1859 <= 32'h0;
    end else begin
      if (11'h743 == _T_12323) begin
        mem_1859 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1860 <= 32'h0;
    end else begin
      if (11'h744 == _T_12323) begin
        mem_1860 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1861 <= 32'h0;
    end else begin
      if (11'h745 == _T_12323) begin
        mem_1861 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1862 <= 32'h0;
    end else begin
      if (11'h746 == _T_12323) begin
        mem_1862 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1863 <= 32'h0;
    end else begin
      if (11'h747 == _T_12323) begin
        mem_1863 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1864 <= 32'h0;
    end else begin
      if (11'h748 == _T_12323) begin
        mem_1864 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1865 <= 32'h0;
    end else begin
      if (11'h749 == _T_12323) begin
        mem_1865 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1866 <= 32'h0;
    end else begin
      if (11'h74a == _T_12323) begin
        mem_1866 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1867 <= 32'h0;
    end else begin
      if (11'h74b == _T_12323) begin
        mem_1867 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1868 <= 32'h0;
    end else begin
      if (11'h74c == _T_12323) begin
        mem_1868 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1869 <= 32'h0;
    end else begin
      if (11'h74d == _T_12323) begin
        mem_1869 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1870 <= 32'h0;
    end else begin
      if (11'h74e == _T_12323) begin
        mem_1870 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1871 <= 32'h0;
    end else begin
      if (11'h74f == _T_12323) begin
        mem_1871 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1872 <= 32'h0;
    end else begin
      if (11'h750 == _T_12323) begin
        mem_1872 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1873 <= 32'h0;
    end else begin
      if (11'h751 == _T_12323) begin
        mem_1873 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1874 <= 32'h0;
    end else begin
      if (11'h752 == _T_12323) begin
        mem_1874 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1875 <= 32'h0;
    end else begin
      if (11'h753 == _T_12323) begin
        mem_1875 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1876 <= 32'h0;
    end else begin
      if (11'h754 == _T_12323) begin
        mem_1876 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1877 <= 32'h0;
    end else begin
      if (11'h755 == _T_12323) begin
        mem_1877 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1878 <= 32'h0;
    end else begin
      if (11'h756 == _T_12323) begin
        mem_1878 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1879 <= 32'h0;
    end else begin
      if (11'h757 == _T_12323) begin
        mem_1879 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1880 <= 32'h0;
    end else begin
      if (11'h758 == _T_12323) begin
        mem_1880 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1881 <= 32'h0;
    end else begin
      if (11'h759 == _T_12323) begin
        mem_1881 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1882 <= 32'h0;
    end else begin
      if (11'h75a == _T_12323) begin
        mem_1882 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1883 <= 32'h0;
    end else begin
      if (11'h75b == _T_12323) begin
        mem_1883 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1884 <= 32'h0;
    end else begin
      if (11'h75c == _T_12323) begin
        mem_1884 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1885 <= 32'h0;
    end else begin
      if (11'h75d == _T_12323) begin
        mem_1885 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1886 <= 32'h0;
    end else begin
      if (11'h75e == _T_12323) begin
        mem_1886 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1887 <= 32'h0;
    end else begin
      if (11'h75f == _T_12323) begin
        mem_1887 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1888 <= 32'h0;
    end else begin
      if (11'h760 == _T_12323) begin
        mem_1888 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1889 <= 32'h0;
    end else begin
      if (11'h761 == _T_12323) begin
        mem_1889 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1890 <= 32'h0;
    end else begin
      if (11'h762 == _T_12323) begin
        mem_1890 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1891 <= 32'h0;
    end else begin
      if (11'h763 == _T_12323) begin
        mem_1891 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1892 <= 32'h0;
    end else begin
      if (11'h764 == _T_12323) begin
        mem_1892 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1893 <= 32'h0;
    end else begin
      if (11'h765 == _T_12323) begin
        mem_1893 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1894 <= 32'h0;
    end else begin
      if (11'h766 == _T_12323) begin
        mem_1894 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1895 <= 32'h0;
    end else begin
      if (11'h767 == _T_12323) begin
        mem_1895 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1896 <= 32'h0;
    end else begin
      if (11'h768 == _T_12323) begin
        mem_1896 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1897 <= 32'h0;
    end else begin
      if (11'h769 == _T_12323) begin
        mem_1897 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1898 <= 32'h0;
    end else begin
      if (11'h76a == _T_12323) begin
        mem_1898 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1899 <= 32'h0;
    end else begin
      if (11'h76b == _T_12323) begin
        mem_1899 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1900 <= 32'h0;
    end else begin
      if (11'h76c == _T_12323) begin
        mem_1900 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1901 <= 32'h0;
    end else begin
      if (11'h76d == _T_12323) begin
        mem_1901 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1902 <= 32'h0;
    end else begin
      if (11'h76e == _T_12323) begin
        mem_1902 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1903 <= 32'h0;
    end else begin
      if (11'h76f == _T_12323) begin
        mem_1903 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1904 <= 32'h0;
    end else begin
      if (11'h770 == _T_12323) begin
        mem_1904 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1905 <= 32'h0;
    end else begin
      if (11'h771 == _T_12323) begin
        mem_1905 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1906 <= 32'h0;
    end else begin
      if (11'h772 == _T_12323) begin
        mem_1906 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1907 <= 32'h0;
    end else begin
      if (11'h773 == _T_12323) begin
        mem_1907 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1908 <= 32'h0;
    end else begin
      if (11'h774 == _T_12323) begin
        mem_1908 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1909 <= 32'h0;
    end else begin
      if (11'h775 == _T_12323) begin
        mem_1909 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1910 <= 32'h0;
    end else begin
      if (11'h776 == _T_12323) begin
        mem_1910 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1911 <= 32'h0;
    end else begin
      if (11'h777 == _T_12323) begin
        mem_1911 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1912 <= 32'h0;
    end else begin
      if (11'h778 == _T_12323) begin
        mem_1912 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1913 <= 32'h0;
    end else begin
      if (11'h779 == _T_12323) begin
        mem_1913 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1914 <= 32'h0;
    end else begin
      if (11'h77a == _T_12323) begin
        mem_1914 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1915 <= 32'h0;
    end else begin
      if (11'h77b == _T_12323) begin
        mem_1915 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1916 <= 32'h0;
    end else begin
      if (11'h77c == _T_12323) begin
        mem_1916 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1917 <= 32'h0;
    end else begin
      if (11'h77d == _T_12323) begin
        mem_1917 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1918 <= 32'h0;
    end else begin
      if (11'h77e == _T_12323) begin
        mem_1918 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1919 <= 32'h0;
    end else begin
      if (11'h77f == _T_12323) begin
        mem_1919 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1920 <= 32'h0;
    end else begin
      if (11'h780 == _T_12323) begin
        mem_1920 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1921 <= 32'h0;
    end else begin
      if (11'h781 == _T_12323) begin
        mem_1921 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1922 <= 32'h0;
    end else begin
      if (11'h782 == _T_12323) begin
        mem_1922 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1923 <= 32'h0;
    end else begin
      if (11'h783 == _T_12323) begin
        mem_1923 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1924 <= 32'h0;
    end else begin
      if (11'h784 == _T_12323) begin
        mem_1924 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1925 <= 32'h0;
    end else begin
      if (11'h785 == _T_12323) begin
        mem_1925 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1926 <= 32'h0;
    end else begin
      if (11'h786 == _T_12323) begin
        mem_1926 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1927 <= 32'h0;
    end else begin
      if (11'h787 == _T_12323) begin
        mem_1927 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1928 <= 32'h0;
    end else begin
      if (11'h788 == _T_12323) begin
        mem_1928 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1929 <= 32'h0;
    end else begin
      if (11'h789 == _T_12323) begin
        mem_1929 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1930 <= 32'h0;
    end else begin
      if (11'h78a == _T_12323) begin
        mem_1930 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1931 <= 32'h0;
    end else begin
      if (11'h78b == _T_12323) begin
        mem_1931 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1932 <= 32'h0;
    end else begin
      if (11'h78c == _T_12323) begin
        mem_1932 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1933 <= 32'h0;
    end else begin
      if (11'h78d == _T_12323) begin
        mem_1933 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1934 <= 32'h0;
    end else begin
      if (11'h78e == _T_12323) begin
        mem_1934 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1935 <= 32'h0;
    end else begin
      if (11'h78f == _T_12323) begin
        mem_1935 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1936 <= 32'h0;
    end else begin
      if (11'h790 == _T_12323) begin
        mem_1936 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1937 <= 32'h0;
    end else begin
      if (11'h791 == _T_12323) begin
        mem_1937 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1938 <= 32'h0;
    end else begin
      if (11'h792 == _T_12323) begin
        mem_1938 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1939 <= 32'h0;
    end else begin
      if (11'h793 == _T_12323) begin
        mem_1939 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1940 <= 32'h0;
    end else begin
      if (11'h794 == _T_12323) begin
        mem_1940 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1941 <= 32'h0;
    end else begin
      if (11'h795 == _T_12323) begin
        mem_1941 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1942 <= 32'h0;
    end else begin
      if (11'h796 == _T_12323) begin
        mem_1942 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1943 <= 32'h0;
    end else begin
      if (11'h797 == _T_12323) begin
        mem_1943 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1944 <= 32'h0;
    end else begin
      if (11'h798 == _T_12323) begin
        mem_1944 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1945 <= 32'h0;
    end else begin
      if (11'h799 == _T_12323) begin
        mem_1945 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1946 <= 32'h0;
    end else begin
      if (11'h79a == _T_12323) begin
        mem_1946 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1947 <= 32'h0;
    end else begin
      if (11'h79b == _T_12323) begin
        mem_1947 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1948 <= 32'h0;
    end else begin
      if (11'h79c == _T_12323) begin
        mem_1948 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1949 <= 32'h0;
    end else begin
      if (11'h79d == _T_12323) begin
        mem_1949 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1950 <= 32'h0;
    end else begin
      if (11'h79e == _T_12323) begin
        mem_1950 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1951 <= 32'h0;
    end else begin
      if (11'h79f == _T_12323) begin
        mem_1951 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1952 <= 32'h0;
    end else begin
      if (11'h7a0 == _T_12323) begin
        mem_1952 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1953 <= 32'h0;
    end else begin
      if (11'h7a1 == _T_12323) begin
        mem_1953 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1954 <= 32'h0;
    end else begin
      if (11'h7a2 == _T_12323) begin
        mem_1954 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1955 <= 32'h0;
    end else begin
      if (11'h7a3 == _T_12323) begin
        mem_1955 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1956 <= 32'h0;
    end else begin
      if (11'h7a4 == _T_12323) begin
        mem_1956 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1957 <= 32'h0;
    end else begin
      if (11'h7a5 == _T_12323) begin
        mem_1957 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1958 <= 32'h0;
    end else begin
      if (11'h7a6 == _T_12323) begin
        mem_1958 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1959 <= 32'h0;
    end else begin
      if (11'h7a7 == _T_12323) begin
        mem_1959 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1960 <= 32'h0;
    end else begin
      if (11'h7a8 == _T_12323) begin
        mem_1960 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1961 <= 32'h0;
    end else begin
      if (11'h7a9 == _T_12323) begin
        mem_1961 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1962 <= 32'h0;
    end else begin
      if (11'h7aa == _T_12323) begin
        mem_1962 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1963 <= 32'h0;
    end else begin
      if (11'h7ab == _T_12323) begin
        mem_1963 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1964 <= 32'h0;
    end else begin
      if (11'h7ac == _T_12323) begin
        mem_1964 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1965 <= 32'h0;
    end else begin
      if (11'h7ad == _T_12323) begin
        mem_1965 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1966 <= 32'h0;
    end else begin
      if (11'h7ae == _T_12323) begin
        mem_1966 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1967 <= 32'h0;
    end else begin
      if (11'h7af == _T_12323) begin
        mem_1967 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1968 <= 32'h0;
    end else begin
      if (11'h7b0 == _T_12323) begin
        mem_1968 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1969 <= 32'h0;
    end else begin
      if (11'h7b1 == _T_12323) begin
        mem_1969 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1970 <= 32'h0;
    end else begin
      if (11'h7b2 == _T_12323) begin
        mem_1970 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1971 <= 32'h0;
    end else begin
      if (11'h7b3 == _T_12323) begin
        mem_1971 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1972 <= 32'h0;
    end else begin
      if (11'h7b4 == _T_12323) begin
        mem_1972 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1973 <= 32'h0;
    end else begin
      if (11'h7b5 == _T_12323) begin
        mem_1973 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1974 <= 32'h0;
    end else begin
      if (11'h7b6 == _T_12323) begin
        mem_1974 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1975 <= 32'h0;
    end else begin
      if (11'h7b7 == _T_12323) begin
        mem_1975 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1976 <= 32'h0;
    end else begin
      if (11'h7b8 == _T_12323) begin
        mem_1976 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1977 <= 32'h0;
    end else begin
      if (11'h7b9 == _T_12323) begin
        mem_1977 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1978 <= 32'h0;
    end else begin
      if (11'h7ba == _T_12323) begin
        mem_1978 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1979 <= 32'h0;
    end else begin
      if (11'h7bb == _T_12323) begin
        mem_1979 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1980 <= 32'h0;
    end else begin
      if (11'h7bc == _T_12323) begin
        mem_1980 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1981 <= 32'h0;
    end else begin
      if (11'h7bd == _T_12323) begin
        mem_1981 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1982 <= 32'h0;
    end else begin
      if (11'h7be == _T_12323) begin
        mem_1982 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1983 <= 32'h0;
    end else begin
      if (11'h7bf == _T_12323) begin
        mem_1983 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1984 <= 32'h0;
    end else begin
      if (11'h7c0 == _T_12323) begin
        mem_1984 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1985 <= 32'h0;
    end else begin
      if (11'h7c1 == _T_12323) begin
        mem_1985 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1986 <= 32'h0;
    end else begin
      if (11'h7c2 == _T_12323) begin
        mem_1986 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1987 <= 32'h0;
    end else begin
      if (11'h7c3 == _T_12323) begin
        mem_1987 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1988 <= 32'h0;
    end else begin
      if (11'h7c4 == _T_12323) begin
        mem_1988 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1989 <= 32'h0;
    end else begin
      if (11'h7c5 == _T_12323) begin
        mem_1989 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1990 <= 32'h0;
    end else begin
      if (11'h7c6 == _T_12323) begin
        mem_1990 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1991 <= 32'h0;
    end else begin
      if (11'h7c7 == _T_12323) begin
        mem_1991 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1992 <= 32'h0;
    end else begin
      if (11'h7c8 == _T_12323) begin
        mem_1992 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1993 <= 32'h0;
    end else begin
      if (11'h7c9 == _T_12323) begin
        mem_1993 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1994 <= 32'h0;
    end else begin
      if (11'h7ca == _T_12323) begin
        mem_1994 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1995 <= 32'h0;
    end else begin
      if (11'h7cb == _T_12323) begin
        mem_1995 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1996 <= 32'h0;
    end else begin
      if (11'h7cc == _T_12323) begin
        mem_1996 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1997 <= 32'h0;
    end else begin
      if (11'h7cd == _T_12323) begin
        mem_1997 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1998 <= 32'h0;
    end else begin
      if (11'h7ce == _T_12323) begin
        mem_1998 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_1999 <= 32'h0;
    end else begin
      if (11'h7cf == _T_12323) begin
        mem_1999 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2000 <= 32'h0;
    end else begin
      if (11'h7d0 == _T_12323) begin
        mem_2000 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2001 <= 32'h0;
    end else begin
      if (11'h7d1 == _T_12323) begin
        mem_2001 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2002 <= 32'h0;
    end else begin
      if (11'h7d2 == _T_12323) begin
        mem_2002 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2003 <= 32'h0;
    end else begin
      if (11'h7d3 == _T_12323) begin
        mem_2003 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2004 <= 32'h0;
    end else begin
      if (11'h7d4 == _T_12323) begin
        mem_2004 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2005 <= 32'h0;
    end else begin
      if (11'h7d5 == _T_12323) begin
        mem_2005 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2006 <= 32'h0;
    end else begin
      if (11'h7d6 == _T_12323) begin
        mem_2006 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2007 <= 32'h0;
    end else begin
      if (11'h7d7 == _T_12323) begin
        mem_2007 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2008 <= 32'h0;
    end else begin
      if (11'h7d8 == _T_12323) begin
        mem_2008 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2009 <= 32'h0;
    end else begin
      if (11'h7d9 == _T_12323) begin
        mem_2009 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2010 <= 32'h0;
    end else begin
      if (11'h7da == _T_12323) begin
        mem_2010 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2011 <= 32'h0;
    end else begin
      if (11'h7db == _T_12323) begin
        mem_2011 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2012 <= 32'h0;
    end else begin
      if (11'h7dc == _T_12323) begin
        mem_2012 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2013 <= 32'h0;
    end else begin
      if (11'h7dd == _T_12323) begin
        mem_2013 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2014 <= 32'h0;
    end else begin
      if (11'h7de == _T_12323) begin
        mem_2014 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2015 <= 32'h0;
    end else begin
      if (11'h7df == _T_12323) begin
        mem_2015 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2016 <= 32'h0;
    end else begin
      if (11'h7e0 == _T_12323) begin
        mem_2016 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2017 <= 32'h0;
    end else begin
      if (11'h7e1 == _T_12323) begin
        mem_2017 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2018 <= 32'h0;
    end else begin
      if (11'h7e2 == _T_12323) begin
        mem_2018 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2019 <= 32'h0;
    end else begin
      if (11'h7e3 == _T_12323) begin
        mem_2019 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2020 <= 32'h0;
    end else begin
      if (11'h7e4 == _T_12323) begin
        mem_2020 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2021 <= 32'h0;
    end else begin
      if (11'h7e5 == _T_12323) begin
        mem_2021 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2022 <= 32'h0;
    end else begin
      if (11'h7e6 == _T_12323) begin
        mem_2022 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2023 <= 32'h0;
    end else begin
      if (11'h7e7 == _T_12323) begin
        mem_2023 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2024 <= 32'h0;
    end else begin
      if (11'h7e8 == _T_12323) begin
        mem_2024 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2025 <= 32'h0;
    end else begin
      if (11'h7e9 == _T_12323) begin
        mem_2025 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2026 <= 32'h0;
    end else begin
      if (11'h7ea == _T_12323) begin
        mem_2026 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2027 <= 32'h0;
    end else begin
      if (11'h7eb == _T_12323) begin
        mem_2027 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2028 <= 32'h0;
    end else begin
      if (11'h7ec == _T_12323) begin
        mem_2028 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2029 <= 32'h0;
    end else begin
      if (11'h7ed == _T_12323) begin
        mem_2029 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2030 <= 32'h0;
    end else begin
      if (11'h7ee == _T_12323) begin
        mem_2030 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2031 <= 32'h0;
    end else begin
      if (11'h7ef == _T_12323) begin
        mem_2031 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2032 <= 32'h0;
    end else begin
      if (11'h7f0 == _T_12323) begin
        mem_2032 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2033 <= 32'h0;
    end else begin
      if (11'h7f1 == _T_12323) begin
        mem_2033 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2034 <= 32'h0;
    end else begin
      if (11'h7f2 == _T_12323) begin
        mem_2034 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2035 <= 32'h0;
    end else begin
      if (11'h7f3 == _T_12323) begin
        mem_2035 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2036 <= 32'h0;
    end else begin
      if (11'h7f4 == _T_12323) begin
        mem_2036 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2037 <= 32'h0;
    end else begin
      if (11'h7f5 == _T_12323) begin
        mem_2037 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2038 <= 32'h0;
    end else begin
      if (11'h7f6 == _T_12323) begin
        mem_2038 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2039 <= 32'h0;
    end else begin
      if (11'h7f7 == _T_12323) begin
        mem_2039 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2040 <= 32'h0;
    end else begin
      if (11'h7f8 == _T_12323) begin
        mem_2040 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2041 <= 32'h0;
    end else begin
      if (11'h7f9 == _T_12323) begin
        mem_2041 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2042 <= 32'h0;
    end else begin
      if (11'h7fa == _T_12323) begin
        mem_2042 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2043 <= 32'h0;
    end else begin
      if (11'h7fb == _T_12323) begin
        mem_2043 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2044 <= 32'h0;
    end else begin
      if (11'h7fc == _T_12323) begin
        mem_2044 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2045 <= 32'h0;
    end else begin
      if (11'h7fd == _T_12323) begin
        mem_2045 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2046 <= 32'h0;
    end else begin
      if (11'h7fe == _T_12323) begin
        mem_2046 <= _GEN_4;
      end
    end
    if (reset) begin
      mem_2047 <= 32'h0;
    end else begin
      if (11'h7ff == _T_12323) begin
        mem_2047 <= _GEN_4;
      end
    end
  end
endmodule
